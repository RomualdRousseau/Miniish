// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     May 30 2022 22:04:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__42118;
    wire N__42117;
    wire N__42116;
    wire N__42107;
    wire N__42106;
    wire N__42105;
    wire N__42098;
    wire N__42097;
    wire N__42096;
    wire N__42089;
    wire N__42088;
    wire N__42087;
    wire N__42080;
    wire N__42079;
    wire N__42078;
    wire N__42071;
    wire N__42070;
    wire N__42069;
    wire N__42062;
    wire N__42061;
    wire N__42060;
    wire N__42053;
    wire N__42052;
    wire N__42051;
    wire N__42044;
    wire N__42043;
    wire N__42042;
    wire N__42035;
    wire N__42034;
    wire N__42033;
    wire N__42026;
    wire N__42025;
    wire N__42024;
    wire N__42017;
    wire N__42016;
    wire N__42015;
    wire N__42008;
    wire N__42007;
    wire N__42006;
    wire N__41999;
    wire N__41998;
    wire N__41997;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41981;
    wire N__41980;
    wire N__41979;
    wire N__41972;
    wire N__41971;
    wire N__41970;
    wire N__41963;
    wire N__41962;
    wire N__41961;
    wire N__41954;
    wire N__41953;
    wire N__41952;
    wire N__41945;
    wire N__41944;
    wire N__41943;
    wire N__41936;
    wire N__41935;
    wire N__41934;
    wire N__41927;
    wire N__41926;
    wire N__41925;
    wire N__41918;
    wire N__41917;
    wire N__41916;
    wire N__41909;
    wire N__41908;
    wire N__41907;
    wire N__41900;
    wire N__41899;
    wire N__41898;
    wire N__41891;
    wire N__41890;
    wire N__41889;
    wire N__41882;
    wire N__41881;
    wire N__41880;
    wire N__41873;
    wire N__41872;
    wire N__41871;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41855;
    wire N__41854;
    wire N__41853;
    wire N__41846;
    wire N__41845;
    wire N__41844;
    wire N__41837;
    wire N__41836;
    wire N__41835;
    wire N__41828;
    wire N__41827;
    wire N__41826;
    wire N__41819;
    wire N__41818;
    wire N__41817;
    wire N__41810;
    wire N__41809;
    wire N__41808;
    wire N__41801;
    wire N__41800;
    wire N__41799;
    wire N__41792;
    wire N__41791;
    wire N__41790;
    wire N__41783;
    wire N__41782;
    wire N__41781;
    wire N__41774;
    wire N__41773;
    wire N__41772;
    wire N__41765;
    wire N__41764;
    wire N__41763;
    wire N__41756;
    wire N__41755;
    wire N__41754;
    wire N__41747;
    wire N__41746;
    wire N__41745;
    wire N__41738;
    wire N__41737;
    wire N__41736;
    wire N__41729;
    wire N__41728;
    wire N__41727;
    wire N__41720;
    wire N__41719;
    wire N__41718;
    wire N__41711;
    wire N__41710;
    wire N__41709;
    wire N__41702;
    wire N__41701;
    wire N__41700;
    wire N__41693;
    wire N__41692;
    wire N__41691;
    wire N__41684;
    wire N__41683;
    wire N__41682;
    wire N__41675;
    wire N__41674;
    wire N__41673;
    wire N__41666;
    wire N__41665;
    wire N__41664;
    wire N__41657;
    wire N__41656;
    wire N__41655;
    wire N__41638;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41626;
    wire N__41623;
    wire N__41620;
    wire N__41617;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41604;
    wire N__41603;
    wire N__41602;
    wire N__41601;
    wire N__41598;
    wire N__41597;
    wire N__41596;
    wire N__41593;
    wire N__41592;
    wire N__41591;
    wire N__41590;
    wire N__41589;
    wire N__41588;
    wire N__41587;
    wire N__41586;
    wire N__41585;
    wire N__41584;
    wire N__41583;
    wire N__41582;
    wire N__41581;
    wire N__41580;
    wire N__41577;
    wire N__41576;
    wire N__41575;
    wire N__41574;
    wire N__41573;
    wire N__41570;
    wire N__41569;
    wire N__41568;
    wire N__41567;
    wire N__41566;
    wire N__41565;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41554;
    wire N__41553;
    wire N__41552;
    wire N__41549;
    wire N__41548;
    wire N__41545;
    wire N__41540;
    wire N__41535;
    wire N__41526;
    wire N__41523;
    wire N__41510;
    wire N__41503;
    wire N__41500;
    wire N__41495;
    wire N__41486;
    wire N__41483;
    wire N__41478;
    wire N__41473;
    wire N__41470;
    wire N__41469;
    wire N__41468;
    wire N__41465;
    wire N__41462;
    wire N__41459;
    wire N__41448;
    wire N__41439;
    wire N__41438;
    wire N__41437;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41419;
    wire N__41414;
    wire N__41407;
    wire N__41402;
    wire N__41399;
    wire N__41398;
    wire N__41395;
    wire N__41390;
    wire N__41385;
    wire N__41382;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41230;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41222;
    wire N__41219;
    wire N__41216;
    wire N__41213;
    wire N__41208;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41163;
    wire N__41158;
    wire N__41155;
    wire N__41152;
    wire N__41149;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41124;
    wire N__41121;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41108;
    wire N__41101;
    wire N__41098;
    wire N__41095;
    wire N__41092;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41065;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41055;
    wire N__41054;
    wire N__41051;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41039;
    wire N__41036;
    wire N__41033;
    wire N__41030;
    wire N__41029;
    wire N__41026;
    wire N__41023;
    wire N__41020;
    wire N__41017;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40984;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40954;
    wire N__40943;
    wire N__40936;
    wire N__40933;
    wire N__40930;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40912;
    wire N__40911;
    wire N__40910;
    wire N__40909;
    wire N__40908;
    wire N__40907;
    wire N__40906;
    wire N__40905;
    wire N__40888;
    wire N__40887;
    wire N__40886;
    wire N__40885;
    wire N__40884;
    wire N__40883;
    wire N__40882;
    wire N__40881;
    wire N__40880;
    wire N__40879;
    wire N__40876;
    wire N__40869;
    wire N__40856;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40848;
    wire N__40847;
    wire N__40846;
    wire N__40845;
    wire N__40844;
    wire N__40843;
    wire N__40840;
    wire N__40837;
    wire N__40836;
    wire N__40831;
    wire N__40828;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40820;
    wire N__40819;
    wire N__40814;
    wire N__40811;
    wire N__40806;
    wire N__40805;
    wire N__40804;
    wire N__40803;
    wire N__40800;
    wire N__40795;
    wire N__40794;
    wire N__40793;
    wire N__40790;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40771;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40752;
    wire N__40739;
    wire N__40726;
    wire N__40725;
    wire N__40724;
    wire N__40723;
    wire N__40722;
    wire N__40721;
    wire N__40720;
    wire N__40719;
    wire N__40718;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40702;
    wire N__40701;
    wire N__40700;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40683;
    wire N__40676;
    wire N__40665;
    wire N__40664;
    wire N__40653;
    wire N__40650;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40627;
    wire N__40624;
    wire N__40621;
    wire N__40618;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40604;
    wire N__40601;
    wire N__40600;
    wire N__40599;
    wire N__40598;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40575;
    wire N__40574;
    wire N__40571;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40527;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40508;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40489;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40465;
    wire N__40464;
    wire N__40463;
    wire N__40462;
    wire N__40461;
    wire N__40460;
    wire N__40459;
    wire N__40458;
    wire N__40457;
    wire N__40456;
    wire N__40455;
    wire N__40454;
    wire N__40453;
    wire N__40452;
    wire N__40451;
    wire N__40450;
    wire N__40449;
    wire N__40448;
    wire N__40447;
    wire N__40446;
    wire N__40445;
    wire N__40444;
    wire N__40443;
    wire N__40442;
    wire N__40441;
    wire N__40440;
    wire N__40439;
    wire N__40438;
    wire N__40437;
    wire N__40436;
    wire N__40435;
    wire N__40434;
    wire N__40433;
    wire N__40432;
    wire N__40431;
    wire N__40430;
    wire N__40429;
    wire N__40428;
    wire N__40427;
    wire N__40426;
    wire N__40425;
    wire N__40424;
    wire N__40423;
    wire N__40422;
    wire N__40421;
    wire N__40420;
    wire N__40419;
    wire N__40418;
    wire N__40417;
    wire N__40416;
    wire N__40415;
    wire N__40414;
    wire N__40413;
    wire N__40412;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40405;
    wire N__40404;
    wire N__40403;
    wire N__40402;
    wire N__40401;
    wire N__40400;
    wire N__40399;
    wire N__40398;
    wire N__40397;
    wire N__40396;
    wire N__40395;
    wire N__40394;
    wire N__40393;
    wire N__40392;
    wire N__40391;
    wire N__40390;
    wire N__40389;
    wire N__40388;
    wire N__40387;
    wire N__40386;
    wire N__40385;
    wire N__40384;
    wire N__40383;
    wire N__40382;
    wire N__40381;
    wire N__40380;
    wire N__40379;
    wire N__40378;
    wire N__40377;
    wire N__40376;
    wire N__40375;
    wire N__40374;
    wire N__40373;
    wire N__40372;
    wire N__40371;
    wire N__40370;
    wire N__40369;
    wire N__40368;
    wire N__40367;
    wire N__40366;
    wire N__40365;
    wire N__40364;
    wire N__40363;
    wire N__40362;
    wire N__40361;
    wire N__40360;
    wire N__40359;
    wire N__40358;
    wire N__40357;
    wire N__40356;
    wire N__40355;
    wire N__40354;
    wire N__40353;
    wire N__40352;
    wire N__40351;
    wire N__40350;
    wire N__40349;
    wire N__40348;
    wire N__40347;
    wire N__40346;
    wire N__40345;
    wire N__40344;
    wire N__40343;
    wire N__40342;
    wire N__40341;
    wire N__40340;
    wire N__40339;
    wire N__40338;
    wire N__40337;
    wire N__40336;
    wire N__40335;
    wire N__40334;
    wire N__40333;
    wire N__40332;
    wire N__40331;
    wire N__40330;
    wire N__40329;
    wire N__40328;
    wire N__40327;
    wire N__40326;
    wire N__40325;
    wire N__40324;
    wire N__40323;
    wire N__40322;
    wire N__40321;
    wire N__40320;
    wire N__40319;
    wire N__40318;
    wire N__40317;
    wire N__40316;
    wire N__40315;
    wire N__40314;
    wire N__40313;
    wire N__40312;
    wire N__40311;
    wire N__40310;
    wire N__40309;
    wire N__40308;
    wire N__40307;
    wire N__40306;
    wire N__40305;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40301;
    wire N__40300;
    wire N__40299;
    wire N__40298;
    wire N__40297;
    wire N__40296;
    wire N__40295;
    wire N__40294;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40290;
    wire N__40289;
    wire N__40288;
    wire N__40287;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39921;
    wire N__39920;
    wire N__39919;
    wire N__39916;
    wire N__39915;
    wire N__39914;
    wire N__39913;
    wire N__39912;
    wire N__39911;
    wire N__39910;
    wire N__39909;
    wire N__39908;
    wire N__39905;
    wire N__39904;
    wire N__39903;
    wire N__39902;
    wire N__39901;
    wire N__39898;
    wire N__39897;
    wire N__39896;
    wire N__39895;
    wire N__39894;
    wire N__39893;
    wire N__39892;
    wire N__39891;
    wire N__39890;
    wire N__39889;
    wire N__39886;
    wire N__39885;
    wire N__39884;
    wire N__39883;
    wire N__39882;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39809;
    wire N__39804;
    wire N__39801;
    wire N__39796;
    wire N__39795;
    wire N__39794;
    wire N__39793;
    wire N__39792;
    wire N__39791;
    wire N__39790;
    wire N__39789;
    wire N__39788;
    wire N__39787;
    wire N__39786;
    wire N__39785;
    wire N__39784;
    wire N__39783;
    wire N__39782;
    wire N__39781;
    wire N__39780;
    wire N__39779;
    wire N__39778;
    wire N__39777;
    wire N__39776;
    wire N__39775;
    wire N__39774;
    wire N__39773;
    wire N__39772;
    wire N__39771;
    wire N__39770;
    wire N__39769;
    wire N__39768;
    wire N__39767;
    wire N__39766;
    wire N__39765;
    wire N__39764;
    wire N__39763;
    wire N__39762;
    wire N__39761;
    wire N__39760;
    wire N__39759;
    wire N__39758;
    wire N__39757;
    wire N__39756;
    wire N__39755;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39703;
    wire N__39700;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39679;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39516;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39498;
    wire N__39497;
    wire N__39494;
    wire N__39491;
    wire N__39488;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39454;
    wire N__39451;
    wire N__39448;
    wire N__39441;
    wire N__39440;
    wire N__39437;
    wire N__39434;
    wire N__39431;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39399;
    wire N__39394;
    wire N__39385;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39377;
    wire N__39376;
    wire N__39375;
    wire N__39374;
    wire N__39373;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39355;
    wire N__39350;
    wire N__39349;
    wire N__39348;
    wire N__39347;
    wire N__39346;
    wire N__39343;
    wire N__39336;
    wire N__39335;
    wire N__39334;
    wire N__39333;
    wire N__39330;
    wire N__39329;
    wire N__39328;
    wire N__39325;
    wire N__39320;
    wire N__39319;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39313;
    wire N__39312;
    wire N__39309;
    wire N__39308;
    wire N__39307;
    wire N__39298;
    wire N__39293;
    wire N__39286;
    wire N__39283;
    wire N__39280;
    wire N__39277;
    wire N__39272;
    wire N__39271;
    wire N__39270;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39247;
    wire N__39244;
    wire N__39241;
    wire N__39238;
    wire N__39231;
    wire N__39224;
    wire N__39221;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39092;
    wire N__39087;
    wire N__39084;
    wire N__39083;
    wire N__39082;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39068;
    wire N__39061;
    wire N__39058;
    wire N__39057;
    wire N__39056;
    wire N__39053;
    wire N__39050;
    wire N__39047;
    wire N__39046;
    wire N__39041;
    wire N__39038;
    wire N__39035;
    wire N__39034;
    wire N__39033;
    wire N__39032;
    wire N__39029;
    wire N__39024;
    wire N__39017;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38938;
    wire N__38937;
    wire N__38936;
    wire N__38935;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38931;
    wire N__38930;
    wire N__38929;
    wire N__38928;
    wire N__38925;
    wire N__38920;
    wire N__38915;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38900;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38812;
    wire N__38809;
    wire N__38806;
    wire N__38803;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38784;
    wire N__38781;
    wire N__38780;
    wire N__38779;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38769;
    wire N__38766;
    wire N__38765;
    wire N__38764;
    wire N__38761;
    wire N__38760;
    wire N__38755;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38722;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38704;
    wire N__38701;
    wire N__38698;
    wire N__38693;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38677;
    wire N__38674;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38575;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38560;
    wire N__38557;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38537;
    wire N__38534;
    wire N__38529;
    wire N__38526;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38501;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38489;
    wire N__38486;
    wire N__38481;
    wire N__38478;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38442;
    wire N__38441;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38431;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38416;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38356;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38341;
    wire N__38340;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38319;
    wire N__38314;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38301;
    wire N__38298;
    wire N__38293;
    wire N__38290;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38245;
    wire N__38244;
    wire N__38239;
    wire N__38236;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38218;
    wire N__38217;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38034;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37984;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37936;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37846;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37810;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37777;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37743;
    wire N__37740;
    wire N__37737;
    wire N__37732;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37704;
    wire N__37701;
    wire N__37700;
    wire N__37697;
    wire N__37694;
    wire N__37691;
    wire N__37688;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37668;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37626;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37584;
    wire N__37583;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37548;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37535;
    wire N__37530;
    wire N__37529;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37500;
    wire N__37497;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37467;
    wire N__37466;
    wire N__37463;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37445;
    wire N__37442;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37391;
    wire N__37384;
    wire N__37383;
    wire N__37380;
    wire N__37379;
    wire N__37376;
    wire N__37375;
    wire N__37374;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37362;
    wire N__37359;
    wire N__37358;
    wire N__37355;
    wire N__37348;
    wire N__37345;
    wire N__37342;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37313;
    wire N__37306;
    wire N__37305;
    wire N__37304;
    wire N__37303;
    wire N__37302;
    wire N__37301;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37261;
    wire N__37260;
    wire N__37255;
    wire N__37252;
    wire N__37249;
    wire N__37244;
    wire N__37241;
    wire N__37238;
    wire N__37233;
    wire N__37230;
    wire N__37225;
    wire N__37216;
    wire N__37213;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37194;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37183;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37165;
    wire N__37162;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37154;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37140;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37125;
    wire N__37120;
    wire N__37115;
    wire N__37112;
    wire N__37111;
    wire N__37108;
    wire N__37103;
    wire N__37100;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37078;
    wire N__37077;
    wire N__37076;
    wire N__37075;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37064;
    wire N__37063;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37040;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36995;
    wire N__36988;
    wire N__36987;
    wire N__36986;
    wire N__36985;
    wire N__36982;
    wire N__36977;
    wire N__36974;
    wire N__36973;
    wire N__36968;
    wire N__36967;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36946;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36919;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36894;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36886;
    wire N__36885;
    wire N__36882;
    wire N__36879;
    wire N__36876;
    wire N__36875;
    wire N__36872;
    wire N__36867;
    wire N__36864;
    wire N__36861;
    wire N__36858;
    wire N__36853;
    wire N__36844;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36832;
    wire N__36831;
    wire N__36830;
    wire N__36829;
    wire N__36826;
    wire N__36821;
    wire N__36818;
    wire N__36811;
    wire N__36810;
    wire N__36807;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36799;
    wire N__36798;
    wire N__36797;
    wire N__36796;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36778;
    wire N__36777;
    wire N__36776;
    wire N__36775;
    wire N__36770;
    wire N__36767;
    wire N__36762;
    wire N__36757;
    wire N__36750;
    wire N__36739;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36731;
    wire N__36728;
    wire N__36727;
    wire N__36726;
    wire N__36723;
    wire N__36722;
    wire N__36721;
    wire N__36718;
    wire N__36715;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36688;
    wire N__36687;
    wire N__36684;
    wire N__36683;
    wire N__36680;
    wire N__36679;
    wire N__36678;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36670;
    wire N__36669;
    wire N__36668;
    wire N__36667;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36653;
    wire N__36648;
    wire N__36643;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36618;
    wire N__36613;
    wire N__36610;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36582;
    wire N__36581;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36568;
    wire N__36563;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36544;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36519;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36487;
    wire N__36486;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36478;
    wire N__36477;
    wire N__36476;
    wire N__36473;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36453;
    wire N__36450;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36436;
    wire N__36433;
    wire N__36430;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36403;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36372;
    wire N__36367;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36309;
    wire N__36308;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36294;
    wire N__36293;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36278;
    wire N__36275;
    wire N__36270;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36191;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36175;
    wire N__36172;
    wire N__36169;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36157;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36037;
    wire N__36034;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35990;
    wire N__35987;
    wire N__35984;
    wire N__35981;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35932;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35924;
    wire N__35923;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35904;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35848;
    wire N__35847;
    wire N__35846;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35836;
    wire N__35833;
    wire N__35832;
    wire N__35827;
    wire N__35826;
    wire N__35825;
    wire N__35824;
    wire N__35821;
    wire N__35820;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35808;
    wire N__35805;
    wire N__35798;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35762;
    wire N__35761;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35751;
    wire N__35750;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35721;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35694;
    wire N__35693;
    wire N__35692;
    wire N__35683;
    wire N__35680;
    wire N__35679;
    wire N__35676;
    wire N__35675;
    wire N__35672;
    wire N__35671;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35640;
    wire N__35635;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35619;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35609;
    wire N__35608;
    wire N__35603;
    wire N__35602;
    wire N__35599;
    wire N__35598;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35569;
    wire N__35564;
    wire N__35563;
    wire N__35560;
    wire N__35553;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35539;
    wire N__35536;
    wire N__35531;
    wire N__35528;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35512;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35504;
    wire N__35499;
    wire N__35498;
    wire N__35495;
    wire N__35492;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35475;
    wire N__35472;
    wire N__35471;
    wire N__35470;
    wire N__35469;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35450;
    wire N__35447;
    wire N__35444;
    wire N__35439;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35420;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35391;
    wire N__35388;
    wire N__35385;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35334;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35292;
    wire N__35287;
    wire N__35284;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35229;
    wire N__35228;
    wire N__35227;
    wire N__35226;
    wire N__35221;
    wire N__35216;
    wire N__35213;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35199;
    wire N__35196;
    wire N__35193;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35178;
    wire N__35175;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35162;
    wire N__35159;
    wire N__35156;
    wire N__35151;
    wire N__35148;
    wire N__35141;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35125;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35117;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35065;
    wire N__35064;
    wire N__35063;
    wire N__35062;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35050;
    wire N__35047;
    wire N__35042;
    wire N__35039;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34977;
    wire N__34976;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34968;
    wire N__34967;
    wire N__34966;
    wire N__34963;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34957;
    wire N__34956;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34941;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34924;
    wire N__34923;
    wire N__34918;
    wire N__34913;
    wire N__34908;
    wire N__34903;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34869;
    wire N__34858;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34843;
    wire N__34840;
    wire N__34839;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34817;
    wire N__34810;
    wire N__34809;
    wire N__34808;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34795;
    wire N__34794;
    wire N__34793;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34748;
    wire N__34745;
    wire N__34742;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34679;
    wire N__34676;
    wire N__34673;
    wire N__34670;
    wire N__34665;
    wire N__34660;
    wire N__34657;
    wire N__34652;
    wire N__34649;
    wire N__34644;
    wire N__34641;
    wire N__34634;
    wire N__34631;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34613;
    wire N__34610;
    wire N__34603;
    wire N__34600;
    wire N__34595;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34560;
    wire N__34559;
    wire N__34558;
    wire N__34555;
    wire N__34554;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34521;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34500;
    wire N__34499;
    wire N__34496;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34488;
    wire N__34485;
    wire N__34484;
    wire N__34475;
    wire N__34472;
    wire N__34469;
    wire N__34466;
    wire N__34463;
    wire N__34460;
    wire N__34457;
    wire N__34454;
    wire N__34449;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34435;
    wire N__34432;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34424;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34393;
    wire N__34392;
    wire N__34387;
    wire N__34386;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34374;
    wire N__34369;
    wire N__34368;
    wire N__34367;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34355;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34344;
    wire N__34343;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34325;
    wire N__34322;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34300;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34287;
    wire N__34286;
    wire N__34283;
    wire N__34280;
    wire N__34277;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34261;
    wire N__34256;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34213;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34154;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34144;
    wire N__34139;
    wire N__34136;
    wire N__34135;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34124;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34110;
    wire N__34107;
    wire N__34096;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34064;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34037;
    wire N__34030;
    wire N__34027;
    wire N__34022;
    wire N__34019;
    wire N__34016;
    wire N__34013;
    wire N__34012;
    wire N__34011;
    wire N__34006;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33994;
    wire N__33993;
    wire N__33990;
    wire N__33989;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33975;
    wire N__33972;
    wire N__33969;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33942;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33903;
    wire N__33898;
    wire N__33895;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33877;
    wire N__33876;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33833;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33814;
    wire N__33809;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33779;
    wire N__33778;
    wire N__33775;
    wire N__33774;
    wire N__33771;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33751;
    wire N__33748;
    wire N__33747;
    wire N__33746;
    wire N__33745;
    wire N__33742;
    wire N__33739;
    wire N__33734;
    wire N__33731;
    wire N__33726;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33705;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33685;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33649;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33518;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33326;
    wire N__33323;
    wire N__33320;
    wire N__33317;
    wire N__33314;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33278;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33247;
    wire N__33244;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33216;
    wire N__33215;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33102;
    wire N__33099;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33050;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33029;
    wire N__33026;
    wire N__33023;
    wire N__33020;
    wire N__33015;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32994;
    wire N__32991;
    wire N__32990;
    wire N__32989;
    wire N__32986;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32963;
    wire N__32960;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32923;
    wire N__32920;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32903;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32860;
    wire N__32857;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32819;
    wire N__32816;
    wire N__32813;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32722;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32704;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32622;
    wire N__32617;
    wire N__32614;
    wire N__32609;
    wire N__32602;
    wire N__32601;
    wire N__32598;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32575;
    wire N__32572;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32521;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32503;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32485;
    wire N__32482;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32464;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32446;
    wire N__32443;
    wire N__32442;
    wire N__32439;
    wire N__32438;
    wire N__32437;
    wire N__32434;
    wire N__32431;
    wire N__32428;
    wire N__32427;
    wire N__32424;
    wire N__32423;
    wire N__32422;
    wire N__32419;
    wire N__32414;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32395;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32370;
    wire N__32365;
    wire N__32362;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32347;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32325;
    wire N__32322;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32310;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32302;
    wire N__32301;
    wire N__32298;
    wire N__32295;
    wire N__32292;
    wire N__32289;
    wire N__32286;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32268;
    wire N__32267;
    wire N__32266;
    wire N__32263;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32257;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32241;
    wire N__32238;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32194;
    wire N__32193;
    wire N__32190;
    wire N__32189;
    wire N__32186;
    wire N__32185;
    wire N__32184;
    wire N__32183;
    wire N__32180;
    wire N__32177;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32165;
    wire N__32162;
    wire N__32159;
    wire N__32152;
    wire N__32149;
    wire N__32142;
    wire N__32137;
    wire N__32136;
    wire N__32133;
    wire N__32132;
    wire N__32129;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32107;
    wire N__32104;
    wire N__32097;
    wire N__32094;
    wire N__32089;
    wire N__32080;
    wire N__32077;
    wire N__32076;
    wire N__32073;
    wire N__32070;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32058;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32041;
    wire N__32038;
    wire N__32035;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32016;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31884;
    wire N__31881;
    wire N__31880;
    wire N__31877;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31863;
    wire N__31862;
    wire N__31853;
    wire N__31850;
    wire N__31847;
    wire N__31844;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31807;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31799;
    wire N__31794;
    wire N__31791;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31781;
    wire N__31776;
    wire N__31771;
    wire N__31768;
    wire N__31767;
    wire N__31766;
    wire N__31759;
    wire N__31758;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31748;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31727;
    wire N__31722;
    wire N__31719;
    wire N__31718;
    wire N__31717;
    wire N__31716;
    wire N__31713;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31678;
    wire N__31677;
    wire N__31674;
    wire N__31673;
    wire N__31670;
    wire N__31669;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31654;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31632;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31621;
    wire N__31618;
    wire N__31617;
    wire N__31610;
    wire N__31607;
    wire N__31604;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31581;
    wire N__31578;
    wire N__31577;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31552;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31529;
    wire N__31522;
    wire N__31519;
    wire N__31516;
    wire N__31513;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31504;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31486;
    wire N__31485;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31460;
    wire N__31459;
    wire N__31454;
    wire N__31451;
    wire N__31448;
    wire N__31447;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31429;
    wire N__31424;
    wire N__31421;
    wire N__31418;
    wire N__31417;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31400;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31388;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31333;
    wire N__31328;
    wire N__31325;
    wire N__31322;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31291;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31279;
    wire N__31278;
    wire N__31277;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31265;
    wire N__31262;
    wire N__31259;
    wire N__31258;
    wire N__31257;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31232;
    wire N__31231;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31219;
    wire N__31214;
    wire N__31211;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31190;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31165;
    wire N__31158;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31069;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31047;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31022;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31010;
    wire N__31009;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30983;
    wire N__30980;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30950;
    wire N__30949;
    wire N__30946;
    wire N__30941;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30907;
    wire N__30900;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30881;
    wire N__30880;
    wire N__30879;
    wire N__30876;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30866;
    wire N__30863;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30840;
    wire N__30839;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30816;
    wire N__30815;
    wire N__30812;
    wire N__30811;
    wire N__30810;
    wire N__30803;
    wire N__30802;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30751;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30688;
    wire N__30683;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30645;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30633;
    wire N__30632;
    wire N__30629;
    wire N__30628;
    wire N__30627;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30611;
    wire N__30608;
    wire N__30605;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30577;
    wire N__30576;
    wire N__30573;
    wire N__30572;
    wire N__30571;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30556;
    wire N__30547;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30539;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30494;
    wire N__30491;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30450;
    wire N__30449;
    wire N__30448;
    wire N__30447;
    wire N__30446;
    wire N__30445;
    wire N__30444;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30427;
    wire N__30418;
    wire N__30417;
    wire N__30416;
    wire N__30415;
    wire N__30414;
    wire N__30413;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30401;
    wire N__30396;
    wire N__30387;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30366;
    wire N__30365;
    wire N__30364;
    wire N__30361;
    wire N__30360;
    wire N__30359;
    wire N__30356;
    wire N__30351;
    wire N__30344;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30330;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30315;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30266;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30219;
    wire N__30218;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30206;
    wire N__30203;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30183;
    wire N__30182;
    wire N__30179;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30168;
    wire N__30165;
    wire N__30164;
    wire N__30163;
    wire N__30160;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30138;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30120;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30102;
    wire N__30099;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30085;
    wire N__30082;
    wire N__30081;
    wire N__30078;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30067;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30046;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30023;
    wire N__30022;
    wire N__30021;
    wire N__30020;
    wire N__30019;
    wire N__30016;
    wire N__30011;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__30000;
    wire N__29999;
    wire N__29998;
    wire N__29995;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29906;
    wire N__29901;
    wire N__29896;
    wire N__29893;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29861;
    wire N__29858;
    wire N__29851;
    wire N__29848;
    wire N__29847;
    wire N__29844;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29834;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29797;
    wire N__29796;
    wire N__29791;
    wire N__29788;
    wire N__29787;
    wire N__29786;
    wire N__29779;
    wire N__29776;
    wire N__29773;
    wire N__29770;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29756;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29737;
    wire N__29734;
    wire N__29731;
    wire N__29730;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29712;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29675;
    wire N__29674;
    wire N__29671;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29650;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29588;
    wire N__29581;
    wire N__29580;
    wire N__29579;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29561;
    wire N__29560;
    wire N__29557;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29520;
    wire N__29519;
    wire N__29518;
    wire N__29515;
    wire N__29514;
    wire N__29511;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29489;
    wire N__29486;
    wire N__29479;
    wire N__29476;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29455;
    wire N__29452;
    wire N__29451;
    wire N__29450;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29444;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29419;
    wire N__29416;
    wire N__29415;
    wire N__29412;
    wire N__29407;
    wire N__29404;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29385;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29338;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29323;
    wire N__29320;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29289;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29229;
    wire N__29226;
    wire N__29225;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29141;
    wire N__29140;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29116;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29095;
    wire N__29090;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29057;
    wire N__29054;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29039;
    wire N__29036;
    wire N__29033;
    wire N__29030;
    wire N__29025;
    wire N__29022;
    wire N__29015;
    wire N__29010;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28956;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28948;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28933;
    wire N__28930;
    wire N__28921;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28899;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28895;
    wire N__28894;
    wire N__28893;
    wire N__28892;
    wire N__28891;
    wire N__28890;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28806;
    wire N__28805;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28764;
    wire N__28763;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28740;
    wire N__28737;
    wire N__28736;
    wire N__28735;
    wire N__28734;
    wire N__28733;
    wire N__28730;
    wire N__28729;
    wire N__28728;
    wire N__28727;
    wire N__28724;
    wire N__28719;
    wire N__28714;
    wire N__28711;
    wire N__28706;
    wire N__28703;
    wire N__28700;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28674;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28658;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28621;
    wire N__28620;
    wire N__28619;
    wire N__28618;
    wire N__28617;
    wire N__28612;
    wire N__28607;
    wire N__28604;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28464;
    wire N__28463;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28438;
    wire N__28437;
    wire N__28436;
    wire N__28435;
    wire N__28434;
    wire N__28433;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28415;
    wire N__28408;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28396;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28384;
    wire N__28381;
    wire N__28380;
    wire N__28379;
    wire N__28376;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28353;
    wire N__28348;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28299;
    wire N__28296;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28286;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28278;
    wire N__28277;
    wire N__28276;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28246;
    wire N__28243;
    wire N__28236;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28196;
    wire N__28195;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28166;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28106;
    wire N__28101;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28067;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27972;
    wire N__27969;
    wire N__27966;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27944;
    wire N__27943;
    wire N__27942;
    wire N__27939;
    wire N__27938;
    wire N__27935;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27897;
    wire N__27894;
    wire N__27893;
    wire N__27892;
    wire N__27889;
    wire N__27888;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27880;
    wire N__27879;
    wire N__27876;
    wire N__27875;
    wire N__27872;
    wire N__27869;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27855;
    wire N__27854;
    wire N__27853;
    wire N__27852;
    wire N__27851;
    wire N__27848;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27781;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27749;
    wire N__27746;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27730;
    wire N__27727;
    wire N__27718;
    wire N__27713;
    wire N__27708;
    wire N__27703;
    wire N__27696;
    wire N__27695;
    wire N__27690;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27670;
    wire N__27667;
    wire N__27666;
    wire N__27663;
    wire N__27662;
    wire N__27659;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27650;
    wire N__27647;
    wire N__27644;
    wire N__27643;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27619;
    wire N__27616;
    wire N__27615;
    wire N__27614;
    wire N__27613;
    wire N__27612;
    wire N__27611;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27539;
    wire N__27536;
    wire N__27533;
    wire N__27530;
    wire N__27525;
    wire N__27522;
    wire N__27517;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27493;
    wire N__27488;
    wire N__27485;
    wire N__27484;
    wire N__27481;
    wire N__27476;
    wire N__27469;
    wire N__27466;
    wire N__27457;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27410;
    wire N__27409;
    wire N__27408;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27393;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27381;
    wire N__27378;
    wire N__27377;
    wire N__27376;
    wire N__27373;
    wire N__27368;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27320;
    wire N__27317;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27307;
    wire N__27304;
    wire N__27297;
    wire N__27292;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27271;
    wire N__27268;
    wire N__27267;
    wire N__27258;
    wire N__27255;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27236;
    wire N__27235;
    wire N__27234;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27223;
    wire N__27222;
    wire N__27221;
    wire N__27218;
    wire N__27215;
    wire N__27214;
    wire N__27213;
    wire N__27210;
    wire N__27209;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27085;
    wire N__27080;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27064;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27041;
    wire N__27036;
    wire N__27029;
    wire N__27026;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26958;
    wire N__26957;
    wire N__26956;
    wire N__26955;
    wire N__26954;
    wire N__26951;
    wire N__26948;
    wire N__26947;
    wire N__26946;
    wire N__26945;
    wire N__26944;
    wire N__26941;
    wire N__26938;
    wire N__26937;
    wire N__26936;
    wire N__26933;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26921;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26899;
    wire N__26898;
    wire N__26897;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26882;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26837;
    wire N__26832;
    wire N__26829;
    wire N__26822;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26805;
    wire N__26800;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26773;
    wire N__26772;
    wire N__26769;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26746;
    wire N__26745;
    wire N__26742;
    wire N__26741;
    wire N__26740;
    wire N__26737;
    wire N__26736;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26727;
    wire N__26726;
    wire N__26725;
    wire N__26722;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26672;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26603;
    wire N__26596;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26580;
    wire N__26577;
    wire N__26576;
    wire N__26573;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26544;
    wire N__26539;
    wire N__26536;
    wire N__26527;
    wire N__26524;
    wire N__26523;
    wire N__26522;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26514;
    wire N__26513;
    wire N__26512;
    wire N__26509;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26482;
    wire N__26479;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26467;
    wire N__26466;
    wire N__26465;
    wire N__26464;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26379;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26357;
    wire N__26348;
    wire N__26341;
    wire N__26340;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26320;
    wire N__26317;
    wire N__26316;
    wire N__26313;
    wire N__26312;
    wire N__26309;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26278;
    wire N__26275;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26262;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26239;
    wire N__26236;
    wire N__26235;
    wire N__26232;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26219;
    wire N__26218;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26146;
    wire N__26143;
    wire N__26138;
    wire N__26135;
    wire N__26132;
    wire N__26129;
    wire N__26126;
    wire N__26121;
    wire N__26118;
    wire N__26113;
    wire N__26108;
    wire N__26105;
    wire N__26100;
    wire N__26091;
    wire N__26090;
    wire N__26085;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26065;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26052;
    wire N__26051;
    wire N__26050;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26042;
    wire N__26041;
    wire N__26040;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26008;
    wire N__26007;
    wire N__26004;
    wire N__26001;
    wire N__26000;
    wire N__25999;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25946;
    wire N__25941;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25912;
    wire N__25905;
    wire N__25898;
    wire N__25895;
    wire N__25890;
    wire N__25889;
    wire N__25884;
    wire N__25881;
    wire N__25876;
    wire N__25873;
    wire N__25870;
    wire N__25869;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25865;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25857;
    wire N__25854;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25844;
    wire N__25843;
    wire N__25842;
    wire N__25841;
    wire N__25840;
    wire N__25837;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25793;
    wire N__25792;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25775;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25736;
    wire N__25733;
    wire N__25728;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25703;
    wire N__25698;
    wire N__25693;
    wire N__25688;
    wire N__25687;
    wire N__25684;
    wire N__25679;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25662;
    wire N__25659;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25641;
    wire N__25640;
    wire N__25639;
    wire N__25638;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25630;
    wire N__25627;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25577;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25487;
    wire N__25484;
    wire N__25479;
    wire N__25476;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25433;
    wire N__25430;
    wire N__25427;
    wire N__25422;
    wire N__25417;
    wire N__25408;
    wire N__25407;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25367;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25296;
    wire N__25295;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25228;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25220;
    wire N__25215;
    wire N__25212;
    wire N__25207;
    wire N__25204;
    wire N__25203;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25179;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25158;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25131;
    wire N__25130;
    wire N__25129;
    wire N__25126;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25108;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25096;
    wire N__25095;
    wire N__25094;
    wire N__25093;
    wire N__25092;
    wire N__25091;
    wire N__25086;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25066;
    wire N__25065;
    wire N__25064;
    wire N__25063;
    wire N__25062;
    wire N__25061;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25039;
    wire N__25038;
    wire N__25035;
    wire N__25034;
    wire N__25031;
    wire N__25028;
    wire N__25025;
    wire N__25018;
    wire N__25015;
    wire N__25014;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25010;
    wire N__25007;
    wire N__25006;
    wire N__25003;
    wire N__24998;
    wire N__24995;
    wire N__24994;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24976;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24956;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24909;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24903;
    wire N__24902;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24898;
    wire N__24889;
    wire N__24886;
    wire N__24877;
    wire N__24876;
    wire N__24875;
    wire N__24874;
    wire N__24873;
    wire N__24870;
    wire N__24865;
    wire N__24862;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24842;
    wire N__24835;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24823;
    wire N__24820;
    wire N__24819;
    wire N__24816;
    wire N__24815;
    wire N__24812;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24793;
    wire N__24790;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24769;
    wire N__24766;
    wire N__24765;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24757;
    wire N__24754;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24730;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24715;
    wire N__24706;
    wire N__24703;
    wire N__24702;
    wire N__24701;
    wire N__24700;
    wire N__24699;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24658;
    wire N__24657;
    wire N__24656;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24645;
    wire N__24644;
    wire N__24643;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24627;
    wire N__24624;
    wire N__24619;
    wire N__24614;
    wire N__24607;
    wire N__24604;
    wire N__24603;
    wire N__24602;
    wire N__24599;
    wire N__24596;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24582;
    wire N__24575;
    wire N__24572;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24548;
    wire N__24541;
    wire N__24540;
    wire N__24537;
    wire N__24532;
    wire N__24531;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24511;
    wire N__24508;
    wire N__24503;
    wire N__24500;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24461;
    wire N__24454;
    wire N__24451;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24442;
    wire N__24441;
    wire N__24438;
    wire N__24433;
    wire N__24428;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24411;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24387;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24357;
    wire N__24356;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24265;
    wire N__24262;
    wire N__24261;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24252;
    wire N__24249;
    wire N__24244;
    wire N__24235;
    wire N__24234;
    wire N__24233;
    wire N__24230;
    wire N__24223;
    wire N__24218;
    wire N__24215;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24158;
    wire N__24155;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24103;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24085;
    wire N__24082;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24066;
    wire N__24063;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24043;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24031;
    wire N__24028;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24009;
    wire N__24006;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23974;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23954;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23938;
    wire N__23933;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23899;
    wire N__23894;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23874;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23857;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23796;
    wire N__23795;
    wire N__23792;
    wire N__23787;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23769;
    wire N__23768;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23760;
    wire N__23759;
    wire N__23756;
    wire N__23755;
    wire N__23754;
    wire N__23753;
    wire N__23752;
    wire N__23751;
    wire N__23750;
    wire N__23749;
    wire N__23736;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23719;
    wire N__23718;
    wire N__23717;
    wire N__23714;
    wire N__23713;
    wire N__23712;
    wire N__23709;
    wire N__23708;
    wire N__23705;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23694;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23677;
    wire N__23676;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23664;
    wire N__23663;
    wire N__23662;
    wire N__23657;
    wire N__23652;
    wire N__23649;
    wire N__23648;
    wire N__23645;
    wire N__23644;
    wire N__23641;
    wire N__23640;
    wire N__23637;
    wire N__23636;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23614;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23597;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23591;
    wire N__23588;
    wire N__23583;
    wire N__23570;
    wire N__23567;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23542;
    wire N__23537;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23523;
    wire N__23522;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23514;
    wire N__23513;
    wire N__23510;
    wire N__23503;
    wire N__23500;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23481;
    wire N__23478;
    wire N__23477;
    wire N__23476;
    wire N__23475;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23447;
    wire N__23446;
    wire N__23445;
    wire N__23442;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23363;
    wire N__23360;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23315;
    wire N__23312;
    wire N__23305;
    wire N__23302;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23280;
    wire N__23273;
    wire N__23268;
    wire N__23263;
    wire N__23258;
    wire N__23251;
    wire N__23248;
    wire N__23239;
    wire N__23234;
    wire N__23231;
    wire N__23224;
    wire N__23221;
    wire N__23220;
    wire N__23219;
    wire N__23216;
    wire N__23211;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23193;
    wire N__23192;
    wire N__23189;
    wire N__23186;
    wire N__23183;
    wire N__23180;
    wire N__23173;
    wire N__23172;
    wire N__23169;
    wire N__23168;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23152;
    wire N__23149;
    wire N__23148;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23133;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23115;
    wire N__23114;
    wire N__23111;
    wire N__23106;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23082;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23070;
    wire N__23069;
    wire N__23066;
    wire N__23061;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23033;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22965;
    wire N__22964;
    wire N__22961;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22926;
    wire N__22923;
    wire N__22918;
    wire N__22915;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22896;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22877;
    wire N__22870;
    wire N__22867;
    wire N__22866;
    wire N__22865;
    wire N__22864;
    wire N__22863;
    wire N__22862;
    wire N__22861;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22853;
    wire N__22844;
    wire N__22835;
    wire N__22828;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22743;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22670;
    wire N__22663;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22629;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22617;
    wire N__22614;
    wire N__22613;
    wire N__22610;
    wire N__22605;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22488;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22413;
    wire N__22410;
    wire N__22409;
    wire N__22406;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22372;
    wire N__22369;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22315;
    wire N__22312;
    wire N__22307;
    wire N__22304;
    wire N__22299;
    wire N__22296;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22216;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22188;
    wire N__22177;
    wire N__22174;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22166;
    wire N__22165;
    wire N__22164;
    wire N__22163;
    wire N__22162;
    wire N__22161;
    wire N__22160;
    wire N__22159;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22136;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22124;
    wire N__22119;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22094;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21910;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21528;
    wire N__21527;
    wire N__21524;
    wire N__21519;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21452;
    wire N__21449;
    wire N__21448;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21429;
    wire N__21428;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21382;
    wire N__21379;
    wire N__21376;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21311;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21274;
    wire N__21269;
    wire N__21264;
    wire N__21261;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21223;
    wire N__21222;
    wire N__21221;
    wire N__21220;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21201;
    wire N__21200;
    wire N__21197;
    wire N__21196;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21175;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21164;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21128;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21089;
    wire N__21084;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21019;
    wire N__21018;
    wire N__21017;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21013;
    wire N__21012;
    wire N__21011;
    wire N__21010;
    wire N__21009;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20909;
    wire N__20906;
    wire N__20893;
    wire N__20884;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20865;
    wire N__20862;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20837;
    wire N__20836;
    wire N__20835;
    wire N__20834;
    wire N__20833;
    wire N__20832;
    wire N__20831;
    wire N__20828;
    wire N__20825;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20689;
    wire N__20684;
    wire N__20679;
    wire N__20674;
    wire N__20671;
    wire N__20664;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20634;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20581;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20557;
    wire N__20554;
    wire N__20553;
    wire N__20552;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20512;
    wire N__20511;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20485;
    wire N__20484;
    wire N__20483;
    wire N__20480;
    wire N__20479;
    wire N__20478;
    wire N__20475;
    wire N__20474;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20444;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20430;
    wire N__20427;
    wire N__20420;
    wire N__20417;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20364;
    wire N__20363;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20355;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20343;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20303;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20274;
    wire N__20269;
    wire N__20266;
    wire N__20263;
    wire N__20262;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20246;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20234;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20218;
    wire N__20215;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20147;
    wire N__20144;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20069;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20065;
    wire N__20064;
    wire N__20063;
    wire N__20058;
    wire N__20057;
    wire N__20048;
    wire N__20043;
    wire N__20038;
    wire N__20031;
    wire N__20030;
    wire N__20029;
    wire N__20026;
    wire N__20025;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20007;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19974;
    wire N__19971;
    wire N__19966;
    wire N__19959;
    wire N__19956;
    wire N__19955;
    wire N__19952;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19912;
    wire N__19909;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19891;
    wire N__19890;
    wire N__19887;
    wire N__19882;
    wire N__19881;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19853;
    wire N__19850;
    wire N__19849;
    wire N__19848;
    wire N__19843;
    wire N__19840;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19808;
    wire N__19795;
    wire N__19794;
    wire N__19793;
    wire N__19790;
    wire N__19785;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19719;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19671;
    wire N__19666;
    wire N__19665;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19620;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19609;
    wire N__19608;
    wire N__19607;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19593;
    wire N__19590;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19586;
    wire N__19585;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19554;
    wire N__19547;
    wire N__19540;
    wire N__19537;
    wire N__19536;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19494;
    wire N__19489;
    wire N__19488;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19455;
    wire N__19450;
    wire N__19449;
    wire N__19446;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19428;
    wire N__19425;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19225;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19162;
    wire N__19159;
    wire N__19158;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19098;
    wire N__19097;
    wire N__19096;
    wire N__19093;
    wire N__19092;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19056;
    wire N__19055;
    wire N__19054;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19015;
    wire N__19014;
    wire N__19013;
    wire N__19010;
    wire N__19009;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__19001;
    wire N__18998;
    wire N__18997;
    wire N__18992;
    wire N__18991;
    wire N__18990;
    wire N__18989;
    wire N__18988;
    wire N__18987;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18954;
    wire N__18937;
    wire N__18936;
    wire N__18933;
    wire N__18932;
    wire N__18929;
    wire N__18928;
    wire N__18925;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18919;
    wire N__18918;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18884;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18849;
    wire N__18848;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18840;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18828;
    wire N__18823;
    wire N__18820;
    wire N__18819;
    wire N__18816;
    wire N__18815;
    wire N__18810;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18791;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18658;
    wire N__18655;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18645;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18637;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18625;
    wire N__18624;
    wire N__18623;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18608;
    wire N__18607;
    wire N__18604;
    wire N__18599;
    wire N__18594;
    wire N__18585;
    wire N__18582;
    wire N__18571;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18563;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18547;
    wire N__18546;
    wire N__18543;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18535;
    wire N__18534;
    wire N__18529;
    wire N__18528;
    wire N__18527;
    wire N__18526;
    wire N__18525;
    wire N__18524;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18494;
    wire N__18491;
    wire N__18488;
    wire N__18481;
    wire N__18478;
    wire N__18473;
    wire N__18470;
    wire N__18463;
    wire N__18448;
    wire N__18445;
    wire N__18444;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18417;
    wire N__18412;
    wire N__18409;
    wire N__18400;
    wire N__18399;
    wire N__18398;
    wire N__18397;
    wire N__18394;
    wire N__18393;
    wire N__18390;
    wire N__18385;
    wire N__18384;
    wire N__18383;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18375;
    wire N__18370;
    wire N__18365;
    wire N__18364;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18345;
    wire N__18334;
    wire N__18331;
    wire N__18330;
    wire N__18329;
    wire N__18326;
    wire N__18325;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18309;
    wire N__18306;
    wire N__18301;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18282;
    wire N__18281;
    wire N__18278;
    wire N__18273;
    wire N__18268;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18260;
    wire N__18255;
    wire N__18252;
    wire N__18251;
    wire N__18248;
    wire N__18243;
    wire N__18238;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18230;
    wire N__18225;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18210;
    wire N__18209;
    wire N__18208;
    wire N__18205;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18191;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18160;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18133;
    wire N__18130;
    wire N__18129;
    wire N__18128;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18093;
    wire N__18086;
    wire N__18079;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18024;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17997;
    wire N__17996;
    wire N__17995;
    wire N__17994;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17962;
    wire N__17961;
    wire N__17960;
    wire N__17957;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17949;
    wire N__17944;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17934;
    wire N__17931;
    wire N__17928;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17912;
    wire N__17909;
    wire N__17902;
    wire N__17901;
    wire N__17898;
    wire N__17897;
    wire N__17894;
    wire N__17893;
    wire N__17892;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17875;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17853;
    wire N__17852;
    wire N__17847;
    wire N__17846;
    wire N__17843;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17814;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17772;
    wire N__17767;
    wire N__17766;
    wire N__17765;
    wire N__17762;
    wire N__17757;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17739;
    wire N__17734;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17719;
    wire N__17716;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17708;
    wire N__17707;
    wire N__17706;
    wire N__17705;
    wire N__17704;
    wire N__17699;
    wire N__17692;
    wire N__17687;
    wire N__17682;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17645;
    wire N__17644;
    wire N__17643;
    wire N__17642;
    wire N__17639;
    wire N__17634;
    wire N__17627;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17599;
    wire N__17598;
    wire N__17597;
    wire N__17596;
    wire N__17595;
    wire N__17594;
    wire N__17591;
    wire N__17590;
    wire N__17587;
    wire N__17586;
    wire N__17585;
    wire N__17584;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17571;
    wire N__17570;
    wire N__17569;
    wire N__17568;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17530;
    wire N__17529;
    wire N__17526;
    wire N__17521;
    wire N__17520;
    wire N__17517;
    wire N__17516;
    wire N__17513;
    wire N__17512;
    wire N__17503;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17475;
    wire N__17472;
    wire N__17467;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17446;
    wire N__17437;
    wire N__17428;
    wire N__17425;
    wire N__17404;
    wire N__17403;
    wire N__17400;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17394;
    wire N__17393;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17389;
    wire N__17386;
    wire N__17381;
    wire N__17380;
    wire N__17379;
    wire N__17376;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17351;
    wire N__17350;
    wire N__17347;
    wire N__17346;
    wire N__17345;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17335;
    wire N__17330;
    wire N__17327;
    wire N__17326;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17314;
    wire N__17311;
    wire N__17306;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17284;
    wire N__17279;
    wire N__17270;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17178;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17002;
    wire N__17001;
    wire N__16998;
    wire N__16997;
    wire N__16994;
    wire N__16993;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16965;
    wire N__16960;
    wire N__16959;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16891;
    wire N__16890;
    wire N__16889;
    wire N__16886;
    wire N__16881;
    wire N__16878;
    wire N__16873;
    wire N__16870;
    wire N__16869;
    wire N__16866;
    wire N__16861;
    wire N__16860;
    wire N__16859;
    wire N__16858;
    wire N__16857;
    wire N__16856;
    wire N__16855;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16846;
    wire N__16843;
    wire N__16842;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16804;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16775;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16756;
    wire N__16753;
    wire N__16746;
    wire N__16743;
    wire N__16738;
    wire N__16733;
    wire N__16728;
    wire N__16723;
    wire N__16708;
    wire N__16707;
    wire N__16706;
    wire N__16705;
    wire N__16704;
    wire N__16703;
    wire N__16702;
    wire N__16699;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16688;
    wire N__16687;
    wire N__16686;
    wire N__16683;
    wire N__16682;
    wire N__16681;
    wire N__16680;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16633;
    wire N__16624;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16594;
    wire N__16593;
    wire N__16592;
    wire N__16591;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16580;
    wire N__16575;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16565;
    wire N__16558;
    wire N__16555;
    wire N__16550;
    wire N__16547;
    wire N__16542;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16515;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16495;
    wire N__16492;
    wire N__16487;
    wire N__16484;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16400;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16387;
    wire N__16382;
    wire N__16381;
    wire N__16380;
    wire N__16379;
    wire N__16378;
    wire N__16377;
    wire N__16376;
    wire N__16373;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16351;
    wire N__16346;
    wire N__16343;
    wire N__16324;
    wire N__16321;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16313;
    wire N__16308;
    wire N__16305;
    wire N__16300;
    wire N__16299;
    wire N__16298;
    wire N__16297;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16293;
    wire N__16292;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16263;
    wire N__16262;
    wire N__16261;
    wire N__16260;
    wire N__16259;
    wire N__16258;
    wire N__16257;
    wire N__16256;
    wire N__16255;
    wire N__16254;
    wire N__16251;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16161;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16154;
    wire N__16151;
    wire N__16148;
    wire N__16145;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16133;
    wire N__16130;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16102;
    wire N__16099;
    wire N__16098;
    wire N__16097;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16075;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16060;
    wire N__16057;
    wire N__16056;
    wire N__16055;
    wire N__16052;
    wire N__16047;
    wire N__16046;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16030;
    wire N__16027;
    wire N__16026;
    wire N__16025;
    wire N__16024;
    wire N__16023;
    wire N__16020;
    wire N__16015;
    wire N__16010;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15918;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15888;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15876;
    wire N__15873;
    wire N__15870;
    wire N__15869;
    wire N__15864;
    wire N__15861;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15838;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15824;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15797;
    wire N__15784;
    wire N__15783;
    wire N__15782;
    wire N__15779;
    wire N__15774;
    wire N__15773;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15765;
    wire N__15764;
    wire N__15763;
    wire N__15762;
    wire N__15761;
    wire N__15758;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15732;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15688;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15674;
    wire N__15673;
    wire N__15672;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15649;
    wire N__15646;
    wire N__15637;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15627;
    wire N__15622;
    wire N__15621;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15565;
    wire N__15558;
    wire N__15551;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15534;
    wire N__15531;
    wire N__15520;
    wire N__15519;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15515;
    wire N__15514;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15480;
    wire N__15477;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15430;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15422;
    wire N__15417;
    wire N__15412;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15369;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15319;
    wire N__15316;
    wire N__15315;
    wire N__15314;
    wire N__15313;
    wire N__15308;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15285;
    wire N__15282;
    wire N__15271;
    wire N__15270;
    wire N__15269;
    wire N__15268;
    wire N__15265;
    wire N__15264;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15260;
    wire N__15257;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15253;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15235;
    wire N__15232;
    wire N__15225;
    wire N__15220;
    wire N__15205;
    wire N__15202;
    wire N__15201;
    wire N__15200;
    wire N__15199;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15185;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15142;
    wire N__15141;
    wire N__15140;
    wire N__15139;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15133;
    wire N__15128;
    wire N__15125;
    wire N__15118;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15012;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14980;
    wire N__14979;
    wire N__14978;
    wire N__14975;
    wire N__14974;
    wire N__14973;
    wire N__14970;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14959;
    wire N__14958;
    wire N__14955;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14930;
    wire N__14927;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14911;
    wire N__14904;
    wire N__14891;
    wire N__14878;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14830;
    wire N__14827;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14814;
    wire N__14813;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14748;
    wire N__14745;
    wire N__14744;
    wire N__14741;
    wire N__14740;
    wire N__14739;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14722;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14706;
    wire N__14705;
    wire N__14700;
    wire N__14697;
    wire N__14696;
    wire N__14695;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14691;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14667;
    wire N__14664;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14592;
    wire N__14591;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14583;
    wire N__14582;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14570;
    wire N__14569;
    wire N__14568;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14552;
    wire N__14549;
    wire N__14544;
    wire N__14537;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14451;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14434;
    wire N__14431;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14405;
    wire N__14402;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14359;
    wire N__14356;
    wire N__14355;
    wire N__14350;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14304;
    wire N__14303;
    wire N__14302;
    wire N__14301;
    wire N__14294;
    wire N__14293;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14285;
    wire N__14284;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14278;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14266;
    wire N__14265;
    wire N__14264;
    wire N__14259;
    wire N__14252;
    wire N__14243;
    wire N__14236;
    wire N__14227;
    wire N__14224;
    wire N__14223;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14204;
    wire N__14201;
    wire N__14194;
    wire N__14191;
    wire N__14190;
    wire N__14189;
    wire N__14184;
    wire N__14181;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14106;
    wire N__14103;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14065;
    wire N__14064;
    wire N__14063;
    wire N__14062;
    wire N__14061;
    wire N__14056;
    wire N__14053;
    wire N__14046;
    wire N__14041;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14000;
    wire N__13993;
    wire N__13992;
    wire N__13991;
    wire N__13990;
    wire N__13987;
    wire N__13986;
    wire N__13985;
    wire N__13984;
    wire N__13977;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13973;
    wire N__13972;
    wire N__13971;
    wire N__13970;
    wire N__13969;
    wire N__13968;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13956;
    wire N__13953;
    wire N__13944;
    wire N__13935;
    wire N__13930;
    wire N__13927;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13899;
    wire N__13898;
    wire N__13893;
    wire N__13892;
    wire N__13891;
    wire N__13888;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13882;
    wire N__13877;
    wire N__13868;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13854;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13794;
    wire N__13793;
    wire N__13792;
    wire N__13791;
    wire N__13788;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13746;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13717;
    wire N__13716;
    wire N__13715;
    wire N__13712;
    wire N__13711;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13707;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13703;
    wire N__13698;
    wire N__13693;
    wire N__13688;
    wire N__13679;
    wire N__13674;
    wire N__13669;
    wire N__13660;
    wire N__13657;
    wire N__13654;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13639;
    wire N__13636;
    wire N__13633;
    wire N__13632;
    wire N__13629;
    wire N__13628;
    wire N__13625;
    wire N__13620;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13554;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13520;
    wire N__13513;
    wire N__13510;
    wire N__13507;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13493;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13450;
    wire N__13447;
    wire N__13446;
    wire N__13445;
    wire N__13442;
    wire N__13437;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13402;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13326;
    wire N__13325;
    wire N__13322;
    wire N__13317;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire VCCG0;
    wire GNDG0;
    wire \this_vga_signals.g1_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.g3_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axb1_cascade_ ;
    wire \this_vga_signals.g2_1_0_cascade_ ;
    wire \this_vga_signals.g2_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ;
    wire \this_vga_signals.g1_0_0_0_cascade_ ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.g2_1 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_cascade_ ;
    wire \this_vga_signals.g3_2 ;
    wire \this_vga_signals.mult1_un75_sum_axb1_3_cascade_ ;
    wire \this_vga_signals.vaddress_m2_1 ;
    wire \this_vga_signals.if_N_9_i ;
    wire \this_vga_signals.if_m1_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axb2_i_0 ;
    wire \this_vga_signals.g2_3 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb1_3_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_2 ;
    wire \this_vga_signals.g1_1_0 ;
    wire \this_vga_signals.g1_4_cascade_ ;
    wire rgb_c_4;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1 ;
    wire \this_vga_signals.vaddress_m2_2 ;
    wire port_clk_c;
    wire \this_vga_signals.g2 ;
    wire \this_vga_signals.g1 ;
    wire \this_vga_signals.N_935_0 ;
    wire port_data_rw_0_i;
    wire \this_vga_signals.g2_2_0 ;
    wire rgb_c_0;
    wire rgb_c_1;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_ ;
    wire \this_vga_signals.g1_0_0_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_ ;
    wire \this_vga_signals.SUM_2_i_i_1_1_3 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_x0 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0 ;
    wire \this_vga_signals.SUM_2_i_i_1_0_3 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_x1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2_mb_sn ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_3 ;
    wire \this_vga_signals.g1_0_0_2_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.g0_0_0_1_0 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_4_cascade_ ;
    wire \this_vga_signals.g2_1_0 ;
    wire \this_vga_signals.g0_4_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0 ;
    wire \this_vga_signals.g0_0_6 ;
    wire \this_vga_signals.g1_0_0_0_0 ;
    wire \this_vga_signals.mult1_un54_sum_ac0_4 ;
    wire \this_vga_signals.g3_0 ;
    wire \this_vga_signals.N_3_2 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.g2_0_0_0 ;
    wire \this_vga_signals.g3_x0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.g3_x1 ;
    wire \this_vga_signals.mult1_un61_sum_axb2_i ;
    wire \this_vga_signals.mult1_un61_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_cascade_ ;
    wire \this_vga_signals.g0_2 ;
    wire \this_vga_signals.mult1_un68_sum_0_3_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_ac0_1 ;
    wire \this_vga_signals.mult1_un47_sum_c3 ;
    wire \this_vga_signals.mult1_un61_sum_c2_0 ;
    wire \this_vga_signals.g3_0_a2_2_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2 ;
    wire \this_vga_signals.g0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0 ;
    wire \this_vga_signals.if_i4_mux_0 ;
    wire \this_vga_signals.vaddress_N_3_i_0_0_cascade_ ;
    wire \this_vga_signals.g2_4_0 ;
    wire \this_vga_signals.g2_0_0 ;
    wire bfn_3_9_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_3_10_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_2_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.N_1_4_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2_2 ;
    wire \this_vga_signals.N_4_3 ;
    wire \this_vga_signals.g1_1_1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_2 ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.g0_0_i_a5_1 ;
    wire \this_vga_signals.N_8 ;
    wire \this_vga_signals.N_6_0_cascade_ ;
    wire \this_vga_signals.g0_1 ;
    wire \this_vga_signals.g3_0_0 ;
    wire \this_vga_signals.g3_1_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_0_2 ;
    wire \this_vga_signals.mult1_un40_sum_axb1_i ;
    wire \this_vga_signals.g0_15 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axb2_0 ;
    wire rgb_c_3;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_1_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb2_i ;
    wire \this_vga_signals.g3_0_1 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_c_0 ;
    wire \this_vga_signals.mult1_un75_sum_ac0_3_d ;
    wire \this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2 ;
    wire \this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_ ;
    wire \this_vga_signals.vaddress_m6_0 ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.mult1_un61_sum_ac0_4 ;
    wire \this_vga_signals.g0_0 ;
    wire \this_vga_signals.g0_0_0_0 ;
    wire \this_vga_signals.g3 ;
    wire \this_vga_signals.g0_0_0_a2_2_0 ;
    wire \this_vga_signals.g0_6_0_a2_3 ;
    wire \this_vga_signals.N_12_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3 ;
    wire \this_vga_signals.g0_1_1 ;
    wire rgb_c_2;
    wire \this_vga_signals.vsync_1_0_a2_3 ;
    wire \this_vga_signals.vsync_1_0_a2_4 ;
    wire this_vga_signals_vsync_1_i;
    wire \this_vga_signals.if_N_6_0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_0_0 ;
    wire \this_vga_signals.vvisibility_i_o2_1_cascade_ ;
    wire \this_vga_signals.vaddress_m2_e_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.N_822_0_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_9_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_7_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_8_repZ0Z1 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_0_0 ;
    wire \this_vga_signals.r_N_4_mux_1_cascade_ ;
    wire \this_vga_signals.N_24_0_1 ;
    wire \this_vga_signals.un2_hsynclt6_0_cascade_ ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire \this_vga_signals.r_N_4_mux_0 ;
    wire \this_vga_signals.N_24_0_0_cascade_ ;
    wire \this_vga_signals.N_4_2_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.g0_0_i_a5_1_0 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.r_N_4_mux_cascade_ ;
    wire \this_vga_signals.N_24_0 ;
    wire \this_vga_signals.r_N_4_mux ;
    wire \this_vga_signals.N_32_0 ;
    wire \this_vga_signals.N_24_0_2_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c2_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_0_0 ;
    wire \this_vga_signals.g0_23_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ;
    wire \this_vga_signals.g0_1_0_0 ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.g0_0_2_0 ;
    wire \this_vga_signals.un2_hsynclt7 ;
    wire this_vga_signals_hsync_1_i;
    wire rgb_c_5;
    wire \this_vga_signals.if_N_8_i_0_cascade_ ;
    wire \this_vga_signals.if_N_9_0_0_cascade_ ;
    wire bfn_5_9_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_5_10_0_;
    wire \this_vga_signals.un4_hsynclto3_0_cascade_ ;
    wire this_vga_signals_un4_lvisibility_1;
    wire this_vga_signals_M_vcounter_q_8;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire \this_vga_signals.N_935_0_g ;
    wire \this_vga_signals.N_1212_g ;
    wire \this_vga_signals.un4_hsynclto7_0 ;
    wire \this_vga_signals.un4_hsynclt9 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire this_vga_signals_M_vcounter_q_7;
    wire \this_vga_signals.g0_0_2 ;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.g0_0_3_0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9 ;
    wire \this_vga_signals.N_935_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire \this_vga_signals.g0_0_0 ;
    wire M_vcounter_q_esr_RNIQJSA2_0_9;
    wire \this_vga_signals.mult1_un82_sum_c3 ;
    wire \this_vga_signals.d_N_11_cascade_ ;
    wire \this_vga_ramdac.m6 ;
    wire \this_vga_ramdac.N_2687_reto ;
    wire \this_vga_ramdac.N_28_i_reto ;
    wire \this_vga_ramdac.m19 ;
    wire \this_vga_ramdac.N_2690_reto ;
    wire \this_vga_signals.mult1_un61_sum_axb1 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_d7lt4 ;
    wire \this_vga_ramdac.N_2691_reto ;
    wire \this_vga_ramdac.m16 ;
    wire \this_vga_ramdac.N_2689_reto ;
    wire \this_vga_signals.N_822_0 ;
    wire \this_vga_signals.M_lcounter_q_3_i_o2_2_1_1 ;
    wire \this_vga_ramdac.N_24_mux ;
    wire M_pcounter_q_ret_1_RNI4VLK7_cascade_;
    wire \this_vga_ramdac.N_2686_reto ;
    wire \this_vga_ramdac.i2_mux ;
    wire M_pcounter_q_ret_1_RNI4VLK7;
    wire \this_vga_ramdac.N_2688_reto ;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_6 ;
    wire \this_vga_signals.g0_6_0_0 ;
    wire M_hcounter_q_esr_RNIU8TO_9;
    wire M_this_vga_signals_address_2;
    wire M_this_vga_signals_address_0;
    wire M_this_vga_signals_address_3;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_0_0 ;
    wire M_this_vga_signals_address_1;
    wire M_this_vga_signals_address_5;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_1;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_3;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_signals.N_2_8_0_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_2_am ;
    wire \this_vga_signals.haddress_1Z0Z_0 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un89_sum_c3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_0 ;
    wire \this_vga_signals.mult1_un61_sum_0_3 ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_2_bm ;
    wire \this_vga_signals.mult1_un75_sum_c2_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.if_N_8_i_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire \this_vga_signals.if_N_9_1 ;
    wire \this_vga_signals.M_pcounter_q_3_1_cascade_ ;
    wire \this_vga_signals.N_3_0 ;
    wire \this_vga_signals.SUM_3_i_0_0 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_signals.mult1_un68_sum_axbxc3_1_0 ;
    wire N_28_0;
    wire \this_vga_signals.M_hcounter_d7lt7_0 ;
    wire \this_vga_signals.M_lcounter_q_3_i_o2_0_1 ;
    wire \this_vga_signals.pixel_clk_i ;
    wire \this_vga_signals.N_83_1_cascade_ ;
    wire \this_vga_signals.N_2_0 ;
    wire \this_vga_signals.M_pcounter_q_i_2_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire \this_vga_signals.M_pcounter_q_0Z0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.N_809_0_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire N_34_0;
    wire port_nmib_1_i;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_9_21_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_9_22_0_;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire \this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ;
    wire this_pixel_clk_M_counter_q_i_1;
    wire M_this_map_ram_write_data_0;
    wire M_this_map_ram_write_data_3;
    wire M_this_map_ram_write_data_4;
    wire dma_0_i;
    wire \this_vga_signals.N_819_0 ;
    wire \this_vga_signals.N_827_0_cascade_ ;
    wire \this_vga_signals.N_826_0 ;
    wire \this_vga_signals.GZ0Z_406 ;
    wire \this_vga_signals.N_83_1 ;
    wire this_pixel_clk_M_counter_q_0;
    wire M_this_map_ram_write_data_1;
    wire M_this_map_ram_write_data_2;
    wire M_this_map_ram_write_data_7;
    wire M_this_map_ram_write_data_5;
    wire M_this_ppu_vram_data_2;
    wire N_825_0;
    wire this_vga_signals_M_lcounter_q_0;
    wire \this_ppu.N_759_0 ;
    wire this_vga_signals_M_lcounter_q_1;
    wire this_vga_signals_M_vcounter_q_9;
    wire \this_ppu.N_5_4_cascade_ ;
    wire \this_ppu.oam_cache.mem_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ;
    wire M_this_map_ram_read_data_0;
    wire M_this_ppu_spr_addr_6;
    wire \this_spr_ram.mem_out_bus4_2 ;
    wire \this_spr_ram.mem_out_bus0_2 ;
    wire M_state_q_RNIQER3C_9;
    wire M_this_ppu_vram_data_1;
    wire M_this_ppu_vram_data_3;
    wire \this_ppu.N_806 ;
    wire M_this_ppu_vram_data_0;
    wire \this_spr_ram.mem_out_bus4_0 ;
    wire \this_spr_ram.mem_out_bus0_0 ;
    wire M_this_map_ram_read_data_2;
    wire M_this_ppu_spr_addr_8;
    wire M_this_map_ram_read_data_1;
    wire M_this_ppu_spr_addr_7;
    wire M_this_map_ram_read_data_3;
    wire M_this_ppu_spr_addr_9;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_spr_addr_10;
    wire \this_ppu.oam_cache.mem_3 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_3 ;
    wire \this_ppu.oam_cache.mem_2 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2 ;
    wire M_this_map_ram_write_data_6;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ;
    wire \this_spr_ram.mem_out_bus7_2 ;
    wire \this_spr_ram.mem_out_bus3_2 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2 ;
    wire M_this_spr_ram_read_data_2;
    wire M_this_spr_ram_read_data_2_cascade_;
    wire \this_spr_ram.mem_out_bus6_2 ;
    wire \this_spr_ram.mem_out_bus2_2 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ;
    wire \this_spr_ram.mem_out_bus7_0 ;
    wire \this_spr_ram.mem_out_bus3_0 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_ ;
    wire M_this_spr_ram_read_data_0;
    wire \this_spr_ram.mem_out_bus7_1 ;
    wire \this_spr_ram.mem_out_bus3_1 ;
    wire \this_spr_ram.mem_out_bus6_0 ;
    wire \this_spr_ram.mem_out_bus2_0 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ;
    wire M_this_spr_ram_read_data_1;
    wire \this_ppu.un1_M_haddress_q_c3_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c6_cascade_ ;
    wire \this_ppu.un1_M_haddress_q_c3 ;
    wire \this_ppu.un1_M_haddress_q_c2 ;
    wire \this_ppu.M_state_qZ0Z_8 ;
    wire \this_spr_ram.mem_out_bus6_3 ;
    wire \this_spr_ram.mem_out_bus2_3 ;
    wire \this_spr_ram.mem_out_bus6_1 ;
    wire \this_spr_ram.mem_out_bus2_1 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1 ;
    wire \this_spr_ram.mem_WE_6 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ;
    wire M_this_spr_ram_read_data_3;
    wire \this_spr_ram.mem_out_bus4_1 ;
    wire \this_spr_ram.mem_out_bus0_1 ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ;
    wire \this_ppu.un1_M_haddress_q_c6 ;
    wire \this_ppu.N_754_0 ;
    wire \this_ppu.M_last_q_RNIGL6V4 ;
    wire \this_spr_ram.mem_WE_8 ;
    wire M_this_map_ram_read_data_6;
    wire \this_spr_ram.mem_radregZ0Z_12 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire M_this_map_ram_read_data_5;
    wire \this_spr_ram.mem_radregZ0Z_11 ;
    wire M_this_state_d_0_sqmuxa;
    wire \this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_ ;
    wire \this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11 ;
    wire bfn_16_22_0_;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1 ;
    wire \this_ppu.un1_M_count_q_1_cry_6_s1 ;
    wire \this_ppu.M_count_q_RNO_0Z0Z_7 ;
    wire \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_2 ;
    wire \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_ ;
    wire \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_4 ;
    wire \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_6 ;
    wire \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ;
    wire \this_ppu.M_count_qZ0Z_3 ;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire \this_spr_ram.mem_out_bus4_3 ;
    wire \this_spr_ram.mem_out_bus0_3 ;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire \this_spr_ram.mem_out_bus7_3 ;
    wire \this_spr_ram.mem_out_bus3_3 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire \this_spr_ram.mem_WE_10 ;
    wire M_this_spr_ram_write_data_2;
    wire \this_ppu.oam_cache.mem_5 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_5 ;
    wire M_this_spr_ram_write_data_1;
    wire N_609;
    wire \this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11 ;
    wire M_this_data_count_qZ0Z_0;
    wire bfn_17_18_0_;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire bfn_17_19_0_;
    wire M_this_data_count_q_cry_8_THRU_CO;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_qZ0Z_10;
    wire M_this_data_count_q_s_10;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_q_cry_10_THRU_CO;
    wire M_this_data_count_q_cry_10;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_q_cry_11_THRU_CO;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_qZ0Z_9;
    wire M_this_data_count_qZ0Z_4;
    wire \this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11 ;
    wire \this_ppu.N_91 ;
    wire \this_ppu.N_760_0_cascade_ ;
    wire \this_ppu.N_762_0 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_ppu.M_last_q ;
    wire \this_ppu.N_5_4 ;
    wire \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ;
    wire \this_ppu.N_268_i_0_0_cascade_ ;
    wire \this_ppu.M_count_qZ0Z_5 ;
    wire M_this_reset_cond_out_0;
    wire \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ;
    wire \this_ppu.N_1323_0_cascade_ ;
    wire \this_ppu.M_count_qZ0Z_1 ;
    wire \this_ppu.M_count_qZ0Z_7 ;
    wire \this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3 ;
    wire M_this_oam_address_qZ0Z_6;
    wire M_this_oam_address_qZ0Z_7;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire port_enb_c;
    wire this_start_data_delay_M_last_q;
    wire M_this_delay_clk_out_0;
    wire N_309_0_cascade_;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_q_cry_5_THRU_CO;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_qZ0Z_7;
    wire M_this_data_count_q_s_13;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_q_s_8;
    wire N_660_i;
    wire M_this_data_count_qZ0Z_8;
    wire N_257;
    wire \this_ppu.M_state_qZ0Z_7 ;
    wire M_this_oam_address_qZ0Z_1;
    wire M_this_oam_address_qZ0Z_0;
    wire N_314_1;
    wire \this_ppu.N_268_i_0_0 ;
    wire \this_ppu.N_1323_0 ;
    wire \this_ppu.M_count_qZ0Z_0 ;
    wire N_611;
    wire M_this_ppu_oam_addr_4;
    wire M_this_data_tmp_qZ0Z_13;
    wire M_this_oam_ram_write_data_13;
    wire M_this_oam_address_qZ0Z_2;
    wire M_this_oam_address_qZ0Z_3;
    wire un1_M_this_oam_address_q_c2;
    wire un1_M_this_oam_address_q_c4;
    wire M_this_oam_address_qZ0Z_5;
    wire un1_M_this_oam_address_q_c4_cascade_;
    wire M_this_oam_address_qZ0Z_4;
    wire un1_M_this_oam_address_q_c6;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_oam_ram_write_data_18;
    wire M_this_data_tmp_qZ0Z_21;
    wire M_this_oam_ram_write_data_21;
    wire M_this_spr_address_qZ0Z_0;
    wire bfn_19_13_0_;
    wire M_this_spr_address_qZ0Z_1;
    wire un1_M_this_spr_address_q_cry_0;
    wire M_this_spr_address_qZ0Z_2;
    wire un1_M_this_spr_address_q_cry_1;
    wire M_this_spr_address_qZ0Z_3;
    wire un1_M_this_spr_address_q_cry_2;
    wire M_this_spr_address_qZ0Z_4;
    wire un1_M_this_spr_address_q_cry_3;
    wire M_this_spr_address_qZ0Z_5;
    wire un1_M_this_spr_address_q_cry_4;
    wire M_this_spr_address_qZ0Z_6;
    wire un1_M_this_spr_address_q_cry_5;
    wire M_this_spr_address_qZ0Z_7;
    wire un1_M_this_spr_address_q_cry_6;
    wire un1_M_this_spr_address_q_cry_7;
    wire M_this_spr_address_qZ0Z_8;
    wire bfn_19_14_0_;
    wire M_this_spr_address_qZ0Z_9;
    wire un1_M_this_spr_address_q_cry_8;
    wire M_this_spr_address_qZ0Z_10;
    wire un1_M_this_spr_address_q_cry_9;
    wire un1_M_this_spr_address_q_cry_10;
    wire un1_M_this_spr_address_q_cry_11;
    wire un1_M_this_spr_address_q_cry_12;
    wire N_1310_0;
    wire bfn_19_17_0_;
    wire M_this_ppu_vram_addr_1;
    wire M_this_scroll_qZ0Z_9;
    wire \this_ppu.un1_M_hoffset_d_cry_0 ;
    wire M_this_ppu_vram_addr_2;
    wire M_this_scroll_qZ0Z_10;
    wire \this_ppu.un1_M_hoffset_d_cry_1 ;
    wire M_this_ppu_vram_addr_3;
    wire M_this_scroll_qZ0Z_11;
    wire \this_ppu.un1_M_hoffset_d_cry_2 ;
    wire M_this_ppu_vram_addr_4;
    wire M_this_scroll_qZ0Z_12;
    wire \this_ppu.un1_M_hoffset_d_cry_3 ;
    wire M_this_scroll_qZ0Z_13;
    wire M_this_ppu_vram_addr_5;
    wire \this_ppu.un1_M_hoffset_d_cry_4 ;
    wire M_this_scroll_qZ0Z_14;
    wire M_this_ppu_vram_addr_6;
    wire \this_ppu.un1_M_hoffset_d_cry_5 ;
    wire \this_ppu.M_haddress_qZ0Z_7 ;
    wire M_this_scroll_qZ0Z_15;
    wire \this_ppu.un1_M_hoffset_d_cry_6 ;
    wire \this_ppu.un1_M_hoffset_d_cry_7 ;
    wire bfn_19_18_0_;
    wire \this_ppu.oam_cache.mem_1 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_1 ;
    wire \this_ppu.N_61_i_cascade_ ;
    wire \this_ppu.N_769_0 ;
    wire \this_ppu.M_state_q_srsts_i_i_o2_4_2 ;
    wire \this_ppu.M_state_qZ0Z_6 ;
    wire \this_ppu.un1_M_state_q_2_0_cascade_ ;
    wire M_this_ppu_oam_addr_5;
    wire \this_ppu.M_oamcurr_qc_0_1 ;
    wire \this_ppu.un1_M_oamcurr_q_2_c5 ;
    wire \this_ppu.M_oamcurr_qZ0Z_6 ;
    wire N_504_g;
    wire \this_ppu.N_17_0 ;
    wire \this_ppu.N_329_0_cascade_ ;
    wire \this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2 ;
    wire \this_ppu.N_21_0 ;
    wire \this_ppu.un1_M_oamcurr_q_2_c3 ;
    wire \this_ppu.N_23_0 ;
    wire \this_ppu.N_329_0 ;
    wire M_this_ppu_oam_addr_0;
    wire M_this_ppu_oam_addr_1;
    wire \this_ppu.un1_M_state_q_2_0 ;
    wire \this_ppu.N_19_0 ;
    wire \this_ppu.un1_M_vaddress_q_c2_cascade_ ;
    wire M_this_data_tmp_qZ0Z_8;
    wire M_this_oam_ram_write_data_8;
    wire M_this_data_tmp_qZ0Z_9;
    wire M_this_oam_ram_write_data_9;
    wire N_1294_0;
    wire M_this_data_tmp_qZ0Z_14;
    wire M_this_oam_ram_write_data_14;
    wire \this_ppu.oam_cache.mem_6 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_6 ;
    wire \this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_ ;
    wire M_this_state_qZ0Z_8;
    wire N_260;
    wire \this_ppu.N_406 ;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12 ;
    wire dma_axb3;
    wire this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_;
    wire dma_0;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10 ;
    wire \this_ppu.N_414_1_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire \this_ppu.N_267 ;
    wire M_this_ppu_vram_addr_0;
    wire M_this_scroll_qZ0Z_8;
    wire bfn_20_19_0_;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_1 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_2 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_3 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_4 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_5 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_6 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_7 ;
    wire bfn_20_20_0_;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_8 ;
    wire \this_ppu.N_242_0 ;
    wire \this_ppu.oam_cache.mem_4 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_4 ;
    wire \this_ppu.M_hoffset_d_0_sqmuxa_7 ;
    wire \this_ppu.M_state_qZ0Z_9 ;
    wire \this_ppu.N_772_0 ;
    wire \this_ppu.N_760_0 ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire \this_ppu.N_799_cascade_ ;
    wire \this_ppu.N_779_0 ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire \this_ppu.N_255 ;
    wire \this_ppu.N_756_0 ;
    wire \this_ppu.un1_M_vaddress_q_c2 ;
    wire \this_ppu.un1_M_vaddress_q_c5 ;
    wire \this_ppu.M_last_q_RNIITCPC ;
    wire bfn_20_24_0_;
    wire \this_ppu.M_oamidx_qZ0Z_1 ;
    wire \this_ppu.un1_M_oamidx_q_cry_0_THRU_CO ;
    wire \this_ppu.un1_M_oamidx_q_cry_0 ;
    wire \this_ppu.un1_M_oamidx_q_cry_1_THRU_CO ;
    wire \this_ppu.un1_M_oamidx_q_cry_1 ;
    wire \this_ppu.un1_M_oamidx_q_cry_2 ;
    wire \this_ppu.M_oamidx_qZ1Z_2 ;
    wire M_this_ppu_oam_addr_3;
    wire \this_ppu.M_oamidx_qZ0Z_3 ;
    wire M_this_ppu_oam_addr_2;
    wire \this_ppu.M_state_q_srsts_0_a3_0_o2_0_6 ;
    wire \this_ppu.N_228_0_i_1_0 ;
    wire \this_ppu.M_oamidx_qZ0Z_0 ;
    wire N_332_0;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_ ;
    wire \this_ppu.N_405 ;
    wire M_this_state_qZ0Z_12;
    wire \this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_ ;
    wire \this_ppu.N_324_0 ;
    wire \this_ppu.N_424_cascade_ ;
    wire \this_ppu.N_449 ;
    wire M_this_state_q_RNI1G0LZ0Z_1;
    wire \this_ppu.N_341_0 ;
    wire \this_ppu.N_934 ;
    wire M_this_state_qZ0Z_5;
    wire M_this_state_qZ0Z_4;
    wire this_ppu_un20_i_a4_0_a2_0_a2_0_2;
    wire N_311_0_cascade_;
    wire M_this_state_q_RNI244K2Z0Z_10;
    wire M_this_state_qZ0Z_10;
    wire M_this_state_q_RNIR71EZ0Z_10;
    wire \this_ppu.hspr_cry_0_c_inv_RNI1203 ;
    wire bfn_21_17_0_;
    wire M_this_ppu_spr_addr_1;
    wire \this_ppu.hspr_cry_0 ;
    wire \this_ppu.hspr_cry_1 ;
    wire M_this_ppu_spr_addr_2;
    wire \this_ppu.M_oam_cache_read_data_i_9 ;
    wire bfn_21_18_0_;
    wire \this_ppu.un1_M_hoffset_q_2_cry_0 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_1 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_2 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_3 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_4 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_5 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_6 ;
    wire \this_ppu.un1_M_hoffset_q_2_cry_7 ;
    wire \this_ppu.M_hoffset_q_i_8 ;
    wire bfn_21_19_0_;
    wire \this_ppu.un1_M_hoffset_q_2_cry_8 ;
    wire \this_ppu.vspr12_0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0 ;
    wire bfn_21_20_0_;
    wire \this_ppu.un1_oam_data_1_cry_0 ;
    wire \this_ppu.un1_oam_data_1_cry_1 ;
    wire \this_ppu.un1_oam_data_1_cry_2 ;
    wire \this_ppu.un1_oam_data_1_cry_3 ;
    wire \this_ppu.un1_oam_data_1_cry_4 ;
    wire \this_ppu.un1_oam_data_1_cry_5 ;
    wire \this_ppu.un1_oam_data_1_cry_6 ;
    wire \this_ppu.un1_oam_data_1_cry_7 ;
    wire bfn_21_21_0_;
    wire \this_ppu.un1_oam_data_1_cry_8 ;
    wire \this_ppu.un1_oam_data_1_cry_8_THRU_CO ;
    wire \this_ppu.vspr_cry_0_c_inv_RNIFK43 ;
    wire bfn_21_22_0_;
    wire M_this_ppu_spr_addr_4;
    wire \this_ppu.vspr_cry_0 ;
    wire \this_ppu.vspr_cry_1 ;
    wire M_this_ppu_spr_addr_5;
    wire \this_ppu.M_oam_cache_read_data_i_17 ;
    wire \this_ppu.oam_cache.mem_17 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_17 ;
    wire M_this_ppu_vram_addr_7;
    wire bfn_21_23_0_;
    wire \this_ppu.M_vaddress_qZ0Z_1 ;
    wire \this_ppu.un1_M_voffset_d_cry_0 ;
    wire \this_ppu.M_vaddress_qZ0Z_2 ;
    wire \this_ppu.un1_M_voffset_d_cry_1 ;
    wire \this_ppu.M_vaddress_qZ0Z_3 ;
    wire \this_ppu.un1_M_voffset_d_cry_2 ;
    wire \this_ppu.M_vaddress_qZ0Z_4 ;
    wire \this_ppu.un1_M_voffset_d_cry_3 ;
    wire \this_ppu.M_vaddress_qZ0Z_5 ;
    wire \this_ppu.un1_M_voffset_d_cry_4 ;
    wire \this_ppu.M_vaddress_qZ0Z_6 ;
    wire \this_ppu.un1_M_voffset_d_cry_5 ;
    wire \this_ppu.M_vaddress_qZ0Z_7 ;
    wire \this_ppu.un1_M_voffset_d_cry_6 ;
    wire \this_ppu.un1_M_voffset_d_cry_7 ;
    wire bfn_21_24_0_;
    wire \this_ppu.N_756_0_0 ;
    wire M_this_data_tmp_qZ0Z_2;
    wire M_this_oam_ram_write_data_2;
    wire M_this_data_tmp_qZ0Z_16;
    wire M_this_oam_ram_write_data_16;
    wire M_this_data_tmp_qZ0Z_5;
    wire M_this_oam_ram_write_data_5;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_oam_ram_write_data_15;
    wire M_this_data_tmp_qZ0Z_19;
    wire M_this_oam_ram_write_data_19;
    wire N_1286_0;
    wire M_this_map_ram_read_data_7;
    wire \this_ppu.N_511 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_ ;
    wire M_this_state_qZ0Z_6;
    wire M_this_state_qZ0Z_7;
    wire this_ppu_un20_i_a4_0_a3_0_a2_1_1;
    wire port_rw_in;
    wire \this_ppu.N_321_0 ;
    wire \this_ppu.N_328_0 ;
    wire M_this_state_qZ0Z_3;
    wire M_this_state_qZ0Z_2;
    wire \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_ ;
    wire \this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0 ;
    wire \this_ppu.N_416 ;
    wire \this_ppu.M_hoffset_q_i_0 ;
    wire bfn_22_18_0_;
    wire \this_ppu.M_hoffset_q_i_1 ;
    wire \this_ppu.un1_M_hoffset_q_cry_0 ;
    wire \this_ppu.M_hoffset_q_i_2 ;
    wire \this_ppu.un1_M_hoffset_q_cry_1 ;
    wire \this_ppu.M_this_ppu_map_addr_i_0 ;
    wire \this_ppu.un1_M_hoffset_q_cry_2 ;
    wire \this_ppu.M_this_ppu_map_addr_i_1 ;
    wire \this_ppu.un1_M_hoffset_q_cry_3 ;
    wire \this_ppu.M_this_ppu_map_addr_i_2 ;
    wire \this_ppu.un1_M_hoffset_q_cry_4 ;
    wire \this_ppu.M_this_ppu_map_addr_i_3 ;
    wire \this_ppu.un1_M_hoffset_q_cry_5 ;
    wire \this_ppu.M_this_ppu_map_addr_i_4 ;
    wire \this_ppu.un1_M_hoffset_q_cry_6 ;
    wire \this_ppu.un1_M_hoffset_q_cry_7 ;
    wire bfn_22_19_0_;
    wire \this_ppu.vspr16_0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_ac0_13_i ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0 ;
    wire \this_ppu.un1_oam_data_1_6 ;
    wire \this_ppu.un1_oam_data_1_8 ;
    wire \this_ppu.un1_oam_data_1_7 ;
    wire \this_ppu.un1_oam_data_1_5 ;
    wire bfn_22_21_0_;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_1 ;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_2 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0 ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_3 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_4 ;
    wire M_this_ppu_map_addr_3;
    wire \this_ppu.read_data_RNI3DGK1_14 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_5 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_6 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_7 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0 ;
    wire \this_ppu.M_hoffset_qZ0Z_8 ;
    wire bfn_22_22_0_;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_8 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO ;
    wire \this_ppu.oam_cache.mem_18 ;
    wire \this_ppu.M_oam_cache_read_data_18 ;
    wire M_this_scroll_qZ0Z_0;
    wire M_this_scroll_qZ0Z_1;
    wire M_this_scroll_qZ0Z_5;
    wire M_this_scroll_qZ0Z_3;
    wire M_this_scroll_qZ0Z_4;
    wire M_this_scroll_qZ0Z_6;
    wire M_this_scroll_qZ0Z_7;
    wire \this_ppu.M_voffset_q_i_0 ;
    wire bfn_22_24_0_;
    wire \this_ppu.M_voffset_qZ0Z_1 ;
    wire \this_ppu.M_voffset_q_i_1 ;
    wire \this_ppu.un1_M_voffset_q_cry_0 ;
    wire \this_ppu.M_voffset_qZ0Z_2 ;
    wire \this_ppu.M_voffset_q_i_2 ;
    wire \this_ppu.un1_M_voffset_q_cry_1 ;
    wire M_this_ppu_map_addr_5;
    wire \this_ppu.M_this_ppu_map_addr_i_5 ;
    wire \this_ppu.un1_M_voffset_q_cry_2 ;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.M_this_ppu_map_addr_i_6 ;
    wire \this_ppu.un1_M_voffset_q_cry_3 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.M_this_ppu_map_addr_i_7 ;
    wire \this_ppu.un1_M_voffset_q_cry_4 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.M_this_ppu_map_addr_i_8 ;
    wire \this_ppu.un1_M_voffset_q_cry_5 ;
    wire M_this_ppu_map_addr_9;
    wire \this_ppu.M_this_ppu_map_addr_i_9 ;
    wire \this_ppu.un1_M_voffset_q_cry_6 ;
    wire \this_ppu.un1_M_voffset_q_cry_7 ;
    wire \this_ppu.M_voffset_qZ0Z_8 ;
    wire \this_ppu.M_voffset_q_i_8 ;
    wire bfn_22_25_0_;
    wire \this_ppu.un1_M_voffset_q_cry_8 ;
    wire \this_ppu.M_state_d14_1 ;
    wire N_433;
    wire N_438;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_oam_ram_write_data_12;
    wire M_this_scroll_qZ0Z_2;
    wire N_1318_0;
    wire M_this_data_tmp_qZ0Z_0;
    wire M_this_oam_ram_write_data_0;
    wire M_this_data_tmp_qZ0Z_1;
    wire M_this_oam_ram_write_data_1;
    wire N_434;
    wire \this_spr_ram.mem_out_bus5_3 ;
    wire \this_spr_ram.mem_out_bus1_3 ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ;
    wire \this_spr_ram.mem_WE_0 ;
    wire \this_ppu.oam_cache.mem_7 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_7 ;
    wire \this_ppu.hspr ;
    wire M_this_ppu_spr_addr_0;
    wire M_this_spr_ram_write_data_0;
    wire \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2 ;
    wire \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3 ;
    wire \this_ppu.N_510 ;
    wire port_address_in_1;
    wire \this_ppu.N_916 ;
    wire \this_ppu.M_state_q_inv_1 ;
    wire \this_ppu.vspr ;
    wire M_this_ppu_spr_addr_3;
    wire \this_ppu.oam_cache.mem_15 ;
    wire \this_ppu.oam_cache.mem_14 ;
    wire M_this_oam_ram_read_data_22;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_22 ;
    wire M_this_oam_ram_read_data_21;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_21 ;
    wire \this_ppu.un1_M_hoffset_q_9 ;
    wire \this_ppu.un1_M_oam_cache_read_data_c7 ;
    wire \this_ppu.un1_M_hoffset_q_10 ;
    wire \this_ppu.un1_M_oam_cache_read_data_c7_cascade_ ;
    wire M_this_ppu_map_addr_4;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0 ;
    wire \this_ppu.oam_cache.mem_12 ;
    wire \this_ppu.M_hoffset_qZ0Z_2 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0 ;
    wire \this_ppu.oam_cache.mem_9 ;
    wire \this_ppu.oam_cache.mem_8 ;
    wire \this_ppu.oam_cache.mem_13 ;
    wire \this_ppu.un1_M_oam_cache_read_data_c4 ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.un1_M_hoffset_q_8 ;
    wire \this_ppu.un1_M_oam_cache_read_data_c4_cascade_ ;
    wire \this_ppu.un1_M_hoffset_q_7 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0 ;
    wire \this_ppu.read_data_RNI80ET_11 ;
    wire M_this_oam_ram_read_data_11;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_11 ;
    wire \this_ppu.oam_cache.mem_11 ;
    wire \this_ppu.un1_M_hoffset_q_6 ;
    wire \this_ppu.M_hoffset_qZ0Z_1 ;
    wire \this_ppu.un1_M_hoffset_q_4 ;
    wire \this_ppu.un1_M_hoffset_q_0 ;
    wire \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0 ;
    wire \this_ppu.un1_oam_data_1_4_c5_0 ;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_23 ;
    wire port_data_c_0;
    wire port_data_c_1;
    wire \this_ppu.oam_cache.mem_16 ;
    wire \this_ppu.M_oam_cache_read_data_16 ;
    wire M_this_data_tmp_qZ0Z_20;
    wire M_this_oam_ram_write_data_20;
    wire M_this_oam_ram_write_data_7;
    wire M_this_data_tmp_qZ0Z_7;
    wire M_this_oam_ram_write_data_3;
    wire M_this_data_tmp_qZ0Z_3;
    wire M_this_oam_ram_write_data_4;
    wire M_this_data_tmp_qZ0Z_4;
    wire N_1302_0;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_oam_ram_write_data_23;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_17 ;
    wire N_440;
    wire N_437;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_oam_ram_write_data_22;
    wire port_data_c_6;
    wire N_439;
    wire \this_spr_ram.mem_WE_2 ;
    wire \this_spr_ram.mem_WE_4 ;
    wire \this_spr_ram.mem_out_bus5_1 ;
    wire \this_spr_ram.mem_out_bus1_1 ;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ;
    wire \this_spr_ram.mem_WE_14 ;
    wire N_260_0;
    wire M_this_spr_address_qZ0Z_13;
    wire M_this_spr_address_qZ0Z_12;
    wire M_this_spr_address_qZ0Z_11;
    wire \this_spr_ram.mem_WE_12 ;
    wire \this_ppu.N_545 ;
    wire M_this_spr_ram_write_data_3;
    wire port_address_in_4;
    wire port_address_in_0;
    wire \this_ppu.N_610 ;
    wire M_this_state_d_0_sqmuxa_2;
    wire led_c_1;
    wire N_608;
    wire M_this_substate_qZ0;
    wire M_this_state_qZ0Z_13;
    wire M_this_state_qZ0Z_11;
    wire M_this_state_qZ0Z_9;
    wire \this_ppu.oam_cache.mem_10 ;
    wire \this_ppu.un1_M_hoffset_q_5 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_18 ;
    wire M_this_state_qZ0Z_1;
    wire port_data_c_7;
    wire M_this_ctrl_flags_qZ0Z_7;
    wire N_312_0;
    wire M_this_ext_address_qZ0Z_0;
    wire bfn_24_21_0_;
    wire M_this_ext_address_qZ0Z_1;
    wire un1_M_this_ext_address_q_cry_0_THRU_CO;
    wire un1_M_this_ext_address_q_cry_0;
    wire M_this_ext_address_qZ0Z_2;
    wire un1_M_this_ext_address_q_cry_1_THRU_CO;
    wire un1_M_this_ext_address_q_cry_1;
    wire M_this_ext_address_qZ0Z_3;
    wire un1_M_this_ext_address_q_cry_2_THRU_CO;
    wire un1_M_this_ext_address_q_cry_2;
    wire un1_M_this_ext_address_q_cry_3;
    wire un1_M_this_ext_address_q_cry_4;
    wire un1_M_this_ext_address_q_cry_5;
    wire un1_M_this_ext_address_q_cry_6;
    wire un1_M_this_ext_address_q_cry_7;
    wire M_this_ext_address_qZ0Z_8;
    wire un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0;
    wire bfn_24_22_0_;
    wire M_this_ext_address_qZ0Z_9;
    wire un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0;
    wire un1_M_this_ext_address_q_cry_8;
    wire un1_M_this_ext_address_q_cry_9;
    wire un1_M_this_ext_address_q_cry_10;
    wire un1_M_this_ext_address_q_cry_11;
    wire un1_M_this_ext_address_q_cry_12;
    wire M_this_ext_address_qZ0Z_14;
    wire un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0;
    wire un1_M_this_ext_address_q_cry_13;
    wire M_this_ext_address_qZ0Z_15;
    wire un1_M_this_ext_address_q_cry_14;
    wire un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_13 ;
    wire M_this_oam_ram_read_data_15;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_15 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_3 ;
    wire M_this_oam_ram_read_data_8;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_8 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_16 ;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_10 ;
    wire M_this_oam_ram_read_data_25;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_25 ;
    wire M_this_oam_ram_read_data_26;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_26 ;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_oam_ram_write_data_10;
    wire M_this_data_tmp_qZ0Z_6;
    wire M_this_oam_ram_write_data_6;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_oam_ram_write_data_11;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_2 ;
    wire \this_ppu.un12lto7Z0Z_4 ;
    wire M_this_oam_ram_read_data_4;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_4 ;
    wire M_this_oam_ram_read_data_5;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_5 ;
    wire M_this_oam_ram_read_data_6;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_6 ;
    wire M_this_oam_ram_read_data_7;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_7 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_1 ;
    wire M_this_oam_ram_read_data_2;
    wire M_this_oam_ram_read_data_1;
    wire M_this_oam_ram_read_data_3;
    wire M_this_oam_ram_read_data_0;
    wire \this_ppu.un12lto7Z0Z_5 ;
    wire M_this_oam_ram_read_data_27;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_27 ;
    wire \this_ppu.un1_oam_data_1_3 ;
    wire M_this_oam_ram_read_data_29;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_29 ;
    wire \this_ppu.un1_oam_data_1_4 ;
    wire M_this_oam_ram_read_data_31;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_31 ;
    wire M_this_oam_ram_read_data_19;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_19 ;
    wire M_this_oam_ram_read_data_20;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_20 ;
    wire M_this_oam_ram_read_data_24;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_24 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.un1_oam_data_1_2 ;
    wire M_this_data_tmp_qZ0Z_17;
    wire M_this_oam_ram_write_data_17;
    wire \this_ppu.un1_oam_data_1_4_c2 ;
    wire M_this_oam_ram_read_data_30;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_30 ;
    wire M_this_oam_ram_read_data_9;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_9 ;
    wire N_435;
    wire M_this_oam_ram_read_data_17;
    wire M_this_oam_ram_read_data_16;
    wire \this_ppu.un1_oam_data_1_1 ;
    wire \this_spr_ram.mem_out_bus5_2 ;
    wire \this_spr_ram.mem_out_bus1_2 ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ;
    wire \this_spr_ram.mem_out_bus5_0 ;
    wire \this_spr_ram.mem_out_bus1_0 ;
    wire \this_spr_ram.mem_radregZ0Z_13 ;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ;
    wire un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0;
    wire port_data_c_2;
    wire M_this_ext_address_qZ0Z_10;
    wire un1_M_this_ext_address_q_cry_3_THRU_CO;
    wire M_this_ext_address_qZ0Z_4;
    wire un1_M_this_ext_address_q_cry_4_THRU_CO;
    wire M_this_ext_address_qZ0Z_5;
    wire un1_M_this_ext_address_q_cry_5_THRU_CO;
    wire M_this_ext_address_qZ0Z_6;
    wire un1_M_this_ext_address_q_cry_6_THRU_CO;
    wire M_this_ext_address_qZ0Z_7;
    wire un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0;
    wire M_this_ext_address_qZ0Z_11;
    wire un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0;
    wire port_data_c_4;
    wire M_this_ext_address_qZ0Z_12;
    wire N_309_0;
    wire N_311_0;
    wire port_data_c_5;
    wire un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0;
    wire M_this_ext_address_qZ0Z_13;
    wire clk_0_c_g;
    wire M_this_reset_cond_out_g_0;
    wire M_this_oam_ram_read_data_12;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_12 ;
    wire port_data_c_3;
    wire M_this_oam_ram_write_data_0_sqmuxa;
    wire N_436;
    wire M_this_oam_ram_read_data_28;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_28 ;
    wire M_this_oam_ram_read_data_14;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_14 ;
    wire port_address_in_2;
    wire port_address_in_3;
    wire port_address_in_6;
    wire port_address_in_5;
    wire \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0 ;
    wire port_address_in_7;
    wire \this_ppu.N_173 ;
    wire _gnd_net_;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__33298,N__33349,N__33397,N__33448,N__33502,N__34306,N__32923,N__35206,N__33004,N__33073}),
            .WADDR({dangling_wire_13,N__19234,N__19267,N__19297,N__19324,N__19351,N__19381,N__19408,N__18685,N__18715,N__18742}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__19645,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__19768,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__19780,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__19657,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__40442),
            .RE(N__23663),
            .WCLKE(N__22177),
            .WCLK(N__40443),
            .WE(N__23667));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__33292,N__33342,N__33391,N__33442,N__33496,N__34297,N__32916,N__35200,N__32998,N__33067}),
            .WADDR({dangling_wire_55,N__19228,N__19261,N__19291,N__19318,N__19345,N__19375,N__19402,N__18679,N__18709,N__18736}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__19759,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__21706,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__19747,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__19636,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__40452),
            .RE(N__23712),
            .WCLKE(N__22159),
            .WCLK(N__40453),
            .WE(N__23713));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__28480,N__25384,N__30196,N__30091,N__28687,N__28753}),
            .WADDR({dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,N__24298,N__24334,N__25195,N__25150,N__25270,N__25312}),
            .MASK({dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .WDATA({N__31939,N__28996,N__25327,N__33664,N__38065,N__38101,N__29074,N__28570,N__36085,N__38089,N__31960,N__36049,N__36067,N__32005,N__33592,N__33610}),
            .RCLKE(),
            .RCLK(N__40462),
            .RE(N__23753),
            .WCLKE(N__39384),
            .WCLK(N__40463),
            .WE(N__23662));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({M_this_oam_ram_read_data_31,M_this_oam_ram_read_data_30,M_this_oam_ram_read_data_29,M_this_oam_ram_read_data_28,M_this_oam_ram_read_data_27,M_this_oam_ram_read_data_26,M_this_oam_ram_read_data_25,M_this_oam_ram_read_data_24,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,N__28474,N__25378,N__30190,N__30085,N__28681,N__28747}),
            .WADDR({dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,N__24292,N__24328,N__25189,N__25144,N__25264,N__25306}),
            .MASK({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .WDATA({N__36349,N__36184,N__33688,N__36340,N__39163,N__39109,N__33580,N__33700,N__35965,N__36322,N__26974,N__35365,N__31924,N__26995,N__38365,N__31978}),
            .RCLKE(),
            .RCLK(N__40464),
            .RE(N__23595),
            .WCLKE(N__39385),
            .WCLK(N__40465),
            .WE(N__23521));
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_0_physical  (
            .RDATA({\this_ppu.oam_cache.mem_15 ,\this_ppu.oam_cache.mem_14 ,\this_ppu.oam_cache.mem_13 ,\this_ppu.oam_cache.mem_12 ,\this_ppu.oam_cache.mem_11 ,\this_ppu.oam_cache.mem_10 ,\this_ppu.oam_cache.mem_9 ,\this_ppu.oam_cache.mem_8 ,\this_ppu.oam_cache.mem_7 ,\this_ppu.oam_cache.mem_6 ,\this_ppu.oam_cache.mem_5 ,\this_ppu.oam_cache.mem_4 ,\this_ppu.oam_cache.mem_3 ,\this_ppu.oam_cache.mem_2 ,\this_ppu.oam_cache.mem_1 ,\this_ppu.oam_cache.mem_0 }),
            .RADDR({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,N__28783,N__28828,N__28597,N__28861}),
            .WADDR({dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,N__30127,N__30229,N__30307,N__29896}),
            .MASK({dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .WDATA({N__37909,N__41356,N__37927,N__39529,N__34990,N__37858,N__39121,N__37882,N__38290,N__38311,N__38332,N__38026,N__37900,N__38056,N__38272,N__38281}),
            .RCLKE(),
            .RCLK(N__40447),
            .RE(N__23719),
            .WCLKE(N__41601),
            .WCLK(N__40448),
            .WE(N__23751));
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,\this_ppu.oam_cache.mem_18 ,\this_ppu.oam_cache.mem_17 ,\this_ppu.oam_cache.mem_16 }),
            .RADDR({dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,N__28777,N__28822,N__28591,N__28855}),
            .WADDR({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__30121,N__30223,N__30301,N__29889}),
            .MASK({dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208}),
            .WDATA({N__38575,N__39148,N__38161,N__41629,N__38194,N__38119,N__38137,N__38455,N__35635,N__34516,N__34444,N__38473,N__38521,N__36535,N__35953,N__37873}),
            .RCLKE(),
            .RCLK(N__40457),
            .RE(N__23752),
            .WCLKE(N__41552),
            .WCLK(N__40458),
            .WE(N__23514));
    defparam \this_spr_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,\this_spr_ram.mem_out_bus0_1 ,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,\this_spr_ram.mem_out_bus0_0 ,dangling_wire_220,dangling_wire_221,dangling_wire_222}),
            .RADDR({N__20779,N__21008,N__21424,N__21175,N__20350,N__31165,N__31388,N__34727,N__30802,N__30995,N__33994}),
            .WADDR({N__27235,N__27409,N__27642,N__27892,N__25618,N__25864,N__26040,N__26297,N__26467,N__26745,N__26945}),
            .MASK({dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238}),
            .WDATA({dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,N__22945,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,N__33863,dangling_wire_250,dangling_wire_251,dangling_wire_252}),
            .RCLKE(),
            .RCLK(N__40434),
            .RE(N__23718),
            .WCLKE(N__36115),
            .WCLK(N__40435),
            .WE(N__23513));
    defparam \this_spr_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,\this_spr_ram.mem_out_bus0_3 ,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,\this_spr_ram.mem_out_bus0_2 ,dangling_wire_264,dangling_wire_265,dangling_wire_266}),
            .RADDR({N__20838,N__21009,N__21423,N__21176,N__20351,N__31190,N__31417,N__34796,N__30750,N__30949,N__33993}),
            .WADDR({N__27213,N__27377,N__27615,N__27887,N__25604,N__25793,N__26039,N__26278,N__26466,N__26731,N__26944}),
            .MASK({dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282}),
            .WDATA({dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__37111,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,N__22733,dangling_wire_294,dangling_wire_295,dangling_wire_296}),
            .RCLKE(),
            .RCLK(N__40417),
            .RE(N__23676),
            .WCLKE(N__36114),
            .WCLK(N__40418),
            .WE(N__23717));
    defparam \this_spr_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,\this_spr_ram.mem_out_bus1_1 ,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,\this_spr_ram.mem_out_bus1_0 ,dangling_wire_308,dangling_wire_309,dangling_wire_310}),
            .RADDR({N__20780,N__21010,N__21425,N__21201,N__20363,N__31219,N__31447,N__34797,N__30787,N__30983,N__33988}),
            .WADDR({N__27186,N__27376,N__27614,N__27875,N__25584,N__25836,N__26000,N__26231,N__26465,N__26725,N__26911}),
            .MASK({dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326}),
            .WDATA({dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,N__22926,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__33844,dangling_wire_338,dangling_wire_339,dangling_wire_340}),
            .RCLKE(),
            .RCLK(N__40396),
            .RE(N__23675),
            .WCLKE(N__37216),
            .WCLK(N__40397),
            .WE(N__23430));
    defparam \this_spr_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,\this_spr_ram.mem_out_bus1_3 ,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,\this_spr_ram.mem_out_bus1_2 ,dangling_wire_352,dangling_wire_353,dangling_wire_354}),
            .RADDR({N__20815,N__21011,N__21426,N__21202,N__20274,N__31245,N__31473,N__34760,N__30815,N__31010,N__33989}),
            .WADDR({N__27176,N__27307,N__27539,N__27855,N__25555,N__25840,N__25999,N__26239,N__26482,N__26726,N__26893}),
            .MASK({dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370}),
            .WDATA({dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,N__37099,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,N__22707,dangling_wire_382,dangling_wire_383,dangling_wire_384}),
            .RCLKE(),
            .RCLK(N__40376),
            .RE(N__23614),
            .WCLKE(N__37212),
            .WCLK(N__40377),
            .WE(N__23674));
    defparam \this_spr_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,\this_spr_ram.mem_out_bus2_1 ,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,\this_spr_ram.mem_out_bus2_0 ,dangling_wire_396,dangling_wire_397,dangling_wire_398}),
            .RADDR({N__20837,N__20992,N__21409,N__21128,N__20262,N__31231,N__31459,N__34785,N__30866,N__31022,N__34011}),
            .WADDR({N__27221,N__27420,N__27650,N__27879,N__25638,N__25873,N__26050,N__26308,N__26521,N__26748,N__26954}),
            .MASK({dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414}),
            .WDATA({dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__22953,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,N__33876,dangling_wire_426,dangling_wire_427,dangling_wire_428}),
            .RCLKE(),
            .RCLK(N__40388),
            .RE(N__23596),
            .WCLKE(N__22768),
            .WCLK(N__40389),
            .WE(N__23597));
    defparam \this_spr_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,\this_spr_ram.mem_out_bus2_3 ,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,\this_spr_ram.mem_out_bus2_2 ,dangling_wire_440,dangling_wire_441,dangling_wire_442}),
            .RADDR({N__20836,N__21018,N__21410,N__21164,N__20234,N__31232,N__31460,N__34809,N__30880,N__31047,N__34072}),
            .WADDR({N__27223,N__27393,N__27629,N__27847,N__25630,N__25869,N__26049,N__26300,N__26522,N__26740,N__26955}),
            .MASK({dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458}),
            .WDATA({dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,N__37154,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,N__22729,dangling_wire_470,dangling_wire_471,dangling_wire_472}),
            .RCLKE(),
            .RCLK(N__40369),
            .RE(N__23525),
            .WCLKE(N__22764),
            .WCLK(N__40370),
            .WE(N__23523));
    defparam \this_spr_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,\this_spr_ram.mem_out_bus3_1 ,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,\this_spr_ram.mem_out_bus3_0 ,dangling_wire_484,dangling_wire_485,dangling_wire_486}),
            .RADDR({N__20835,N__21019,N__21439,N__21171,N__20302,N__31257,N__31485,N__34810,N__30881,N__31069,N__34087}),
            .WADDR({N__27222,N__27421,N__27651,N__27851,N__25619,N__25868,N__26051,N__26261,N__26513,N__26736,N__26946}),
            .MASK({dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502}),
            .WDATA({dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,N__22964,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,N__33894,dangling_wire_514,dangling_wire_515,dangling_wire_516}),
            .RCLKE(),
            .RCLK(N__40342),
            .RE(N__23524),
            .WCLKE(N__22368),
            .WCLK(N__40343),
            .WE(N__23522));
    defparam \this_spr_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,\this_spr_ram.mem_out_bus3_3 ,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,\this_spr_ram.mem_out_bus3_2 ,dangling_wire_528,dangling_wire_529,dangling_wire_530}),
            .RADDR({N__20805,N__21029,N__21440,N__21200,N__20335,N__31258,N__31486,N__34799,N__30888,N__31086,N__34088}),
            .WADDR({N__27236,N__27438,N__27612,N__27852,N__25641,N__25857,N__26052,N__26312,N__26514,N__26671,N__26947}),
            .MASK({dangling_wire_531,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546}),
            .WDATA({dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,N__37161,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,N__22744,dangling_wire_558,dangling_wire_559,dangling_wire_560}),
            .RCLKE(),
            .RCLK(N__40325),
            .RE(N__23456),
            .WCLKE(N__22372),
            .WCLK(N__40324),
            .WE(N__23447));
    defparam \this_spr_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,\this_spr_ram.mem_out_bus4_1 ,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,\this_spr_ram.mem_out_bus4_0 ,dangling_wire_572,dangling_wire_573,dangling_wire_574}),
            .RADDR({N__20834,N__21030,N__21452,N__21196,N__20355,N__31277,N__31503,N__34800,N__30889,N__31087,N__34095}),
            .WADDR({N__27243,N__27449,N__27662,N__27853,N__25639,N__25853,N__26061,N__26316,N__26523,N__26735,N__26958}),
            .MASK({dangling_wire_575,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590}),
            .WDATA({dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,N__22969,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,N__33898,dangling_wire_602,dangling_wire_603,dangling_wire_604}),
            .RCLKE(),
            .RCLK(N__40310),
            .RE(N__23455),
            .WCLKE(N__22020),
            .WCLK(N__40311),
            .WE(N__23446));
    defparam \this_spr_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,\this_spr_ram.mem_out_bus4_3 ,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,\this_spr_ram.mem_out_bus4_2 ,dangling_wire_616,dangling_wire_617,dangling_wire_618}),
            .RADDR({N__20833,N__21034,N__21453,N__21220,N__20364,N__31278,N__31504,N__34798,N__30839,N__31009,N__34096}),
            .WADDR({N__27247,N__27454,N__27667,N__27854,N__25645,N__25792,N__26062,N__26317,N__26524,N__26747,N__26959}),
            .MASK({dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634}),
            .WDATA({dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,N__37165,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,N__22735,dangling_wire_646,dangling_wire_647,dangling_wire_648}),
            .RCLKE(),
            .RCLK(N__40302),
            .RE(N__23445),
            .WCLKE(N__22024),
            .WCLK(N__40303),
            .WE(N__23363));
    defparam \this_spr_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,\this_spr_ram.mem_out_bus5_1 ,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,\this_spr_ram.mem_out_bus5_0 ,dangling_wire_660,dangling_wire_661,dangling_wire_662}),
            .RADDR({N__20841,N__21012,N__21427,N__21221,N__20312,N__31265,N__31400,N__34795,N__30816,N__31035,N__34012}),
            .WADDR({N__27194,N__27381,N__27619,N__27868,N__25577,N__25841,N__26007,N__26218,N__26456,N__26730,N__26897}),
            .MASK({dangling_wire_663,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678}),
            .WDATA({dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,N__22946,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,N__33864,dangling_wire_690,dangling_wire_691,dangling_wire_692}),
            .RCLKE(),
            .RCLK(N__40351),
            .RE(N__23613),
            .WCLKE(N__36156),
            .WCLK(N__40352),
            .WE(N__23429));
    defparam \this_spr_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,\this_spr_ram.mem_out_bus5_3 ,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,\this_spr_ram.mem_out_bus5_2 ,dangling_wire_704,dangling_wire_705,dangling_wire_706}),
            .RADDR({N__20842,N__21013,N__21428,N__21222,N__20342,N__31279,N__31493,N__34794,N__30840,N__31057,N__34037}),
            .WADDR({N__27214,N__27410,N__27611,N__27880,N__25597,N__25842,N__26008,N__26274,N__26508,N__26672,N__26898}),
            .MASK({dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722}),
            .WDATA({dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,N__37125,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,N__22743,dangling_wire_734,dangling_wire_735,dangling_wire_736}),
            .RCLKE(),
            .RCLK(N__40332),
            .RE(N__23548),
            .WCLKE(N__36157),
            .WCLK(N__40331),
            .WE(N__23546));
    defparam \this_spr_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,\this_spr_ram.mem_out_bus6_1 ,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,\this_spr_ram.mem_out_bus6_0 ,dangling_wire_748,dangling_wire_749,dangling_wire_750}),
            .RADDR({N__20839,N__21014,N__21429,N__21235,N__20346,N__31291,N__31429,N__34808,N__30810,N__31076,N__34064}),
            .WADDR({N__27209,N__27431,N__27643,N__27888,N__25614,N__25865,N__26041,N__26307,N__26489,N__26746,N__26936}),
            .MASK({dangling_wire_751,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766}),
            .WDATA({dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,N__22960,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,N__33877,dangling_wire_778,dangling_wire_779,dangling_wire_780}),
            .RCLKE(),
            .RCLK(N__40319),
            .RE(N__23547),
            .WCLKE(N__36168),
            .WCLK(N__40320),
            .WE(N__23428));
    defparam \this_spr_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,\this_spr_ram.mem_out_bus6_3 ,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,\this_spr_ram.mem_out_bus6_2 ,dangling_wire_792,dangling_wire_793,dangling_wire_794}),
            .RADDR({N__20840,N__21015,N__21447,N__21236,N__20362,N__31301,N__31505,N__34792,N__30811,N__31088,N__34065}),
            .WADDR({N__27234,N__27445,N__27658,N__27893,N__25626,N__25866,N__26042,N__26299,N__26463,N__26749,N__26937}),
            .MASK({dangling_wire_795,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810}),
            .WDATA({dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,N__37140,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,N__22734,dangling_wire_822,dangling_wire_823,dangling_wire_824}),
            .RCLKE(),
            .RCLK(N__40306),
            .RE(N__23476),
            .WCLKE(N__36172),
            .WCLK(N__40307),
            .WE(N__23481));
    defparam \this_spr_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,\this_spr_ram.mem_out_bus7_1 ,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,\this_spr_ram.mem_out_bus7_0 ,dangling_wire_836,dangling_wire_837,dangling_wire_838}),
            .RADDR({N__20831,N__21016,N__21448,N__21243,N__20365,N__31308,N__31512,N__34793,N__30862,N__31095,N__34085}),
            .WADDR({N__27193,N__27453,N__27666,N__27897,N__25637,N__25843,N__26059,N__26235,N__26512,N__26741,N__26956}),
            .MASK({dangling_wire_839,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854}),
            .WDATA({dangling_wire_855,dangling_wire_856,dangling_wire_857,dangling_wire_858,N__22968,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,N__33887,dangling_wire_866,dangling_wire_867,dangling_wire_868}),
            .RCLKE(),
            .RCLK(N__40298),
            .RE(N__23477),
            .WCLKE(N__34213),
            .WCLK(N__40299),
            .WE(N__23405));
    defparam \this_spr_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,\this_spr_ram.mem_out_bus7_3 ,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,\this_spr_ram.mem_out_bus7_2 ,dangling_wire_880,dangling_wire_881,dangling_wire_882}),
            .RADDR({N__20832,N__21017,N__21454,N__21244,N__20325,N__31309,N__31513,N__34807,N__30879,N__31096,N__34086}),
            .WADDR({N__27233,N__27408,N__27613,N__27898,N__25640,N__25867,N__26060,N__26298,N__26464,N__26721,N__26957}),
            .MASK({dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898}),
            .WDATA({dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,N__37153,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,N__22742,dangling_wire_910,dangling_wire_911,dangling_wire_912}),
            .RCLKE(),
            .RCLK(N__40288),
            .RE(N__23545),
            .WCLKE(N__34212),
            .WCLK(N__40289),
            .WE(N__23591));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917,dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,dangling_wire_922,dangling_wire_923,dangling_wire_924,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_925,dangling_wire_926,dangling_wire_927,N__14839,N__18778,N__18013,N__17188,N__17197,N__17215,N__17164,N__17206}),
            .WADDR({dangling_wire_928,dangling_wire_929,dangling_wire_930,N__31863,N__28087,N__28138,N__28213,N__28303,N__28381,N__27961,N__29356}),
            .MASK({dangling_wire_931,dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,dangling_wire_943,dangling_wire_944,dangling_wire_945,dangling_wire_946}),
            .WDATA({dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,N__21544,N__19735,N__20092,N__21514}),
            .RCLKE(),
            .RCLK(N__40293),
            .RE(N__23475),
            .WCLKE(N__20107),
            .WCLK(N__40294),
            .WE(N__23454));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__42116),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__42118),
            .DIN(N__42117),
            .DOUT(N__42116),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__42118),
            .PADOUT(N__42117),
            .PADIN(N__42116),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__42107),
            .DIN(N__42106),
            .DOUT(N__42105),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__42107),
            .PADOUT(N__42106),
            .PADIN(N__42105),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__42098),
            .DIN(N__42097),
            .DOUT(N__42096),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__42098),
            .PADOUT(N__42097),
            .PADIN(N__42096),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__42089),
            .DIN(N__42088),
            .DOUT(N__42087),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__42089),
            .PADOUT(N__42088),
            .PADIN(N__42087),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__17236),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__42080),
            .DIN(N__42079),
            .DOUT(N__42078),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__42080),
            .PADOUT(N__42079),
            .PADIN(N__42078),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15973),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__42071),
            .DIN(N__42070),
            .DOUT(N__42069),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__42071),
            .PADOUT(N__42070),
            .PADIN(N__42069),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__23636),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__42062),
            .DIN(N__42061),
            .DOUT(N__42060),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__42062),
            .PADOUT(N__42061),
            .PADIN(N__42060),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36904),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__42053),
            .DIN(N__42052),
            .DOUT(N__42051),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__42053),
            .PADOUT(N__42052),
            .PADIN(N__42051),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__42044),
            .DIN(N__42043),
            .DOUT(N__42042),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__42044),
            .PADOUT(N__42043),
            .PADIN(N__42042),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__42035),
            .DIN(N__42034),
            .DOUT(N__42033),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__42035),
            .PADOUT(N__42034),
            .PADIN(N__42033),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__42026),
            .DIN(N__42025),
            .DOUT(N__42024),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__42026),
            .PADOUT(N__42025),
            .PADIN(N__42024),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__42017),
            .DIN(N__42016),
            .DOUT(N__42015),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__42017),
            .PADOUT(N__42016),
            .PADIN(N__42015),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__42008),
            .DIN(N__42007),
            .DOUT(N__42006),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__42008),
            .PADOUT(N__42007),
            .PADIN(N__42006),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__41999),
            .DIN(N__41998),
            .DOUT(N__41997),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__41999),
            .PADOUT(N__41998),
            .PADIN(N__41997),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__37717),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19593));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__41990),
            .DIN(N__41989),
            .DOUT(N__41988),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__41990),
            .PADOUT(N__41989),
            .PADIN(N__41988),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__37681),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19620));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__41981),
            .DIN(N__41980),
            .DOUT(N__41979),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__41981),
            .PADOUT(N__41980),
            .PADIN(N__41979),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__37636),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19609));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__41972),
            .DIN(N__41971),
            .DOUT(N__41970),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__41972),
            .PADOUT(N__41971),
            .PADIN(N__41970),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__37600),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19607));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__41963),
            .DIN(N__41962),
            .DOUT(N__41961),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__41963),
            .PADOUT(N__41962),
            .PADIN(N__41961),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__38626),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19588));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__41954),
            .DIN(N__41953),
            .DOUT(N__41952),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__41954),
            .PADOUT(N__41953),
            .PADIN(N__41952),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__41233),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19536));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__41945),
            .DIN(N__41944),
            .DOUT(N__41943),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__41945),
            .PADOUT(N__41944),
            .PADIN(N__41943),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__41191),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19587));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__41936),
            .DIN(N__41935),
            .DOUT(N__41934),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__41936),
            .PADOUT(N__41935),
            .PADIN(N__41934),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__41146),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19585));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__41927),
            .DIN(N__41926),
            .DOUT(N__41925),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__41927),
            .PADOUT(N__41926),
            .PADIN(N__41925),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__38665),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19608));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__41918),
            .DIN(N__41917),
            .DOUT(N__41916),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__41918),
            .PADOUT(N__41917),
            .PADIN(N__41916),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__41092),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19624));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__41909),
            .DIN(N__41908),
            .DOUT(N__41907),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__41909),
            .PADOUT(N__41908),
            .PADIN(N__41907),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40936),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19589));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__41900),
            .DIN(N__41899),
            .DOUT(N__41898),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__41900),
            .PADOUT(N__41899),
            .PADIN(N__41898),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__40492),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19564));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__41891),
            .DIN(N__41890),
            .DOUT(N__41889),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__41891),
            .PADOUT(N__41890),
            .PADIN(N__41889),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__38011),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19586));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__41882),
            .DIN(N__41881),
            .DOUT(N__41880),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__41882),
            .PADOUT(N__41881),
            .PADIN(N__41880),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37975),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19554));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__41873),
            .DIN(N__41872),
            .DOUT(N__41871),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__41873),
            .PADOUT(N__41872),
            .PADIN(N__41871),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37837),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19521));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__41864),
            .DIN(N__41863),
            .DOUT(N__41862),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__41864),
            .PADOUT(N__41863),
            .PADIN(N__41862),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37801),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19619));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__41855),
            .DIN(N__41854),
            .DOUT(N__41853),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__41855),
            .PADOUT(N__41854),
            .PADIN(N__41853),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__41846),
            .DIN(N__41845),
            .DOUT(N__41844),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__41846),
            .PADOUT(N__41845),
            .PADIN(N__41844),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__41837),
            .DIN(N__41836),
            .DOUT(N__41835),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__41837),
            .PADOUT(N__41836),
            .PADIN(N__41835),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__41828),
            .DIN(N__41827),
            .DOUT(N__41826),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__41828),
            .PADOUT(N__41827),
            .PADIN(N__41826),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__41819),
            .DIN(N__41818),
            .DOUT(N__41817),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__41819),
            .PADOUT(N__41818),
            .PADIN(N__41817),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__41810),
            .DIN(N__41809),
            .DOUT(N__41808),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__41810),
            .PADOUT(N__41809),
            .PADIN(N__41808),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__41801),
            .DIN(N__41800),
            .DOUT(N__41799),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__41801),
            .PADOUT(N__41800),
            .PADIN(N__41799),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__41792),
            .DIN(N__41791),
            .DOUT(N__41790),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__41792),
            .PADOUT(N__41791),
            .PADIN(N__41790),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__41783),
            .DIN(N__41782),
            .DOUT(N__41781),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__41783),
            .PADOUT(N__41782),
            .PADIN(N__41781),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__41774),
            .DIN(N__41773),
            .DOUT(N__41772),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__41774),
            .PADOUT(N__41773),
            .PADIN(N__41772),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13423),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__41765),
            .DIN(N__41764),
            .DOUT(N__41763),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__41765),
            .PADOUT(N__41764),
            .PADIN(N__41763),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29239),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__41756),
            .DIN(N__41755),
            .DOUT(N__41754),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__41756),
            .PADOUT(N__41755),
            .PADIN(N__41754),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__41747),
            .DIN(N__41746),
            .DOUT(N__41745),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__41747),
            .PADOUT(N__41746),
            .PADIN(N__41745),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__18760),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__41738),
            .DIN(N__41737),
            .DOUT(N__41736),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__41738),
            .PADOUT(N__41737),
            .PADIN(N__41736),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__23750),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__19488));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__41729),
            .DIN(N__41728),
            .DOUT(N__41727),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__41729),
            .PADOUT(N__41728),
            .PADIN(N__41727),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13399),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__41720),
            .DIN(N__41719),
            .DOUT(N__41718),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__41720),
            .PADOUT(N__41719),
            .PADIN(N__41718),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13387),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__41711),
            .DIN(N__41710),
            .DOUT(N__41709),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__41711),
            .PADOUT(N__41710),
            .PADIN(N__41709),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15094),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__41702),
            .DIN(N__41701),
            .DOUT(N__41700),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__41702),
            .PADOUT(N__41701),
            .PADIN(N__41700),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15031),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__41693),
            .DIN(N__41692),
            .DOUT(N__41691),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__41693),
            .PADOUT(N__41692),
            .PADIN(N__41691),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__13342),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__41684),
            .DIN(N__41683),
            .DOUT(N__41682),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__41684),
            .PADOUT(N__41683),
            .PADIN(N__41682),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15955),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__41675),
            .DIN(N__41674),
            .DOUT(N__41673),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__41675),
            .PADOUT(N__41674),
            .PADIN(N__41673),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__41666),
            .DIN(N__41665),
            .DOUT(N__41664),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__41666),
            .PADOUT(N__41665),
            .PADIN(N__41664),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__16441),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__41657),
            .DIN(N__41656),
            .DOUT(N__41655),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__41657),
            .PADOUT(N__41656),
            .PADIN(N__41655),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__15064),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__10490 (
            .O(N__41638),
            .I(N__41635));
    LocalMux I__10489 (
            .O(N__41635),
            .I(N__41632));
    Odrv4 I__10488 (
            .O(N__41632),
            .I(M_this_oam_ram_read_data_28));
    InMux I__10487 (
            .O(N__41629),
            .I(N__41626));
    LocalMux I__10486 (
            .O(N__41626),
            .I(N__41623));
    Span4Mux_h I__10485 (
            .O(N__41623),
            .I(N__41620));
    Odrv4 I__10484 (
            .O(N__41620),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_28 ));
    InMux I__10483 (
            .O(N__41617),
            .I(N__41614));
    LocalMux I__10482 (
            .O(N__41614),
            .I(N__41611));
    Span4Mux_v I__10481 (
            .O(N__41611),
            .I(N__41608));
    Odrv4 I__10480 (
            .O(N__41608),
            .I(M_this_oam_ram_read_data_14));
    InMux I__10479 (
            .O(N__41605),
            .I(N__41598));
    InMux I__10478 (
            .O(N__41604),
            .I(N__41593));
    CascadeMux I__10477 (
            .O(N__41603),
            .I(N__41577));
    InMux I__10476 (
            .O(N__41602),
            .I(N__41570));
    CEMux I__10475 (
            .O(N__41601),
            .I(N__41561));
    LocalMux I__10474 (
            .O(N__41598),
            .I(N__41558));
    InMux I__10473 (
            .O(N__41597),
            .I(N__41555));
    CascadeMux I__10472 (
            .O(N__41596),
            .I(N__41549));
    LocalMux I__10471 (
            .O(N__41593),
            .I(N__41545));
    InMux I__10470 (
            .O(N__41592),
            .I(N__41540));
    InMux I__10469 (
            .O(N__41591),
            .I(N__41540));
    InMux I__10468 (
            .O(N__41590),
            .I(N__41535));
    InMux I__10467 (
            .O(N__41589),
            .I(N__41535));
    InMux I__10466 (
            .O(N__41588),
            .I(N__41526));
    InMux I__10465 (
            .O(N__41587),
            .I(N__41526));
    InMux I__10464 (
            .O(N__41586),
            .I(N__41526));
    InMux I__10463 (
            .O(N__41585),
            .I(N__41526));
    InMux I__10462 (
            .O(N__41584),
            .I(N__41523));
    InMux I__10461 (
            .O(N__41583),
            .I(N__41510));
    InMux I__10460 (
            .O(N__41582),
            .I(N__41510));
    InMux I__10459 (
            .O(N__41581),
            .I(N__41510));
    InMux I__10458 (
            .O(N__41580),
            .I(N__41510));
    InMux I__10457 (
            .O(N__41577),
            .I(N__41510));
    InMux I__10456 (
            .O(N__41576),
            .I(N__41510));
    InMux I__10455 (
            .O(N__41575),
            .I(N__41503));
    InMux I__10454 (
            .O(N__41574),
            .I(N__41503));
    InMux I__10453 (
            .O(N__41573),
            .I(N__41503));
    LocalMux I__10452 (
            .O(N__41570),
            .I(N__41500));
    InMux I__10451 (
            .O(N__41569),
            .I(N__41495));
    InMux I__10450 (
            .O(N__41568),
            .I(N__41495));
    InMux I__10449 (
            .O(N__41567),
            .I(N__41486));
    InMux I__10448 (
            .O(N__41566),
            .I(N__41486));
    InMux I__10447 (
            .O(N__41565),
            .I(N__41486));
    InMux I__10446 (
            .O(N__41564),
            .I(N__41486));
    LocalMux I__10445 (
            .O(N__41561),
            .I(N__41483));
    Span4Mux_v I__10444 (
            .O(N__41558),
            .I(N__41478));
    LocalMux I__10443 (
            .O(N__41555),
            .I(N__41478));
    InMux I__10442 (
            .O(N__41554),
            .I(N__41473));
    InMux I__10441 (
            .O(N__41553),
            .I(N__41473));
    CEMux I__10440 (
            .O(N__41552),
            .I(N__41470));
    InMux I__10439 (
            .O(N__41549),
            .I(N__41465));
    InMux I__10438 (
            .O(N__41548),
            .I(N__41462));
    Span4Mux_h I__10437 (
            .O(N__41545),
            .I(N__41459));
    LocalMux I__10436 (
            .O(N__41540),
            .I(N__41448));
    LocalMux I__10435 (
            .O(N__41535),
            .I(N__41448));
    LocalMux I__10434 (
            .O(N__41526),
            .I(N__41448));
    LocalMux I__10433 (
            .O(N__41523),
            .I(N__41448));
    LocalMux I__10432 (
            .O(N__41510),
            .I(N__41448));
    LocalMux I__10431 (
            .O(N__41503),
            .I(N__41439));
    Span4Mux_v I__10430 (
            .O(N__41500),
            .I(N__41439));
    LocalMux I__10429 (
            .O(N__41495),
            .I(N__41439));
    LocalMux I__10428 (
            .O(N__41486),
            .I(N__41439));
    Span4Mux_h I__10427 (
            .O(N__41483),
            .I(N__41433));
    Span4Mux_v I__10426 (
            .O(N__41478),
            .I(N__41430));
    LocalMux I__10425 (
            .O(N__41473),
            .I(N__41427));
    LocalMux I__10424 (
            .O(N__41470),
            .I(N__41424));
    InMux I__10423 (
            .O(N__41469),
            .I(N__41419));
    InMux I__10422 (
            .O(N__41468),
            .I(N__41419));
    LocalMux I__10421 (
            .O(N__41465),
            .I(N__41414));
    LocalMux I__10420 (
            .O(N__41462),
            .I(N__41414));
    Span4Mux_h I__10419 (
            .O(N__41459),
            .I(N__41407));
    Span4Mux_v I__10418 (
            .O(N__41448),
            .I(N__41407));
    Span4Mux_v I__10417 (
            .O(N__41439),
            .I(N__41407));
    InMux I__10416 (
            .O(N__41438),
            .I(N__41402));
    InMux I__10415 (
            .O(N__41437),
            .I(N__41402));
    InMux I__10414 (
            .O(N__41436),
            .I(N__41399));
    Span4Mux_h I__10413 (
            .O(N__41433),
            .I(N__41395));
    Span4Mux_h I__10412 (
            .O(N__41430),
            .I(N__41390));
    Span4Mux_v I__10411 (
            .O(N__41427),
            .I(N__41390));
    Span12Mux_s11_v I__10410 (
            .O(N__41424),
            .I(N__41385));
    LocalMux I__10409 (
            .O(N__41419),
            .I(N__41385));
    Span4Mux_v I__10408 (
            .O(N__41414),
            .I(N__41382));
    Span4Mux_h I__10407 (
            .O(N__41407),
            .I(N__41377));
    LocalMux I__10406 (
            .O(N__41402),
            .I(N__41377));
    LocalMux I__10405 (
            .O(N__41399),
            .I(N__41374));
    InMux I__10404 (
            .O(N__41398),
            .I(N__41371));
    Odrv4 I__10403 (
            .O(N__41395),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__10402 (
            .O(N__41390),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv12 I__10401 (
            .O(N__41385),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__10400 (
            .O(N__41382),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__10399 (
            .O(N__41377),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__10398 (
            .O(N__41374),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__10397 (
            .O(N__41371),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    InMux I__10396 (
            .O(N__41356),
            .I(N__41353));
    LocalMux I__10395 (
            .O(N__41353),
            .I(N__41350));
    Span4Mux_h I__10394 (
            .O(N__41350),
            .I(N__41347));
    Odrv4 I__10393 (
            .O(N__41347),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_14 ));
    InMux I__10392 (
            .O(N__41344),
            .I(N__41341));
    LocalMux I__10391 (
            .O(N__41341),
            .I(N__41338));
    Span4Mux_v I__10390 (
            .O(N__41338),
            .I(N__41335));
    Sp12to4 I__10389 (
            .O(N__41335),
            .I(N__41332));
    Span12Mux_s10_h I__10388 (
            .O(N__41332),
            .I(N__41329));
    Odrv12 I__10387 (
            .O(N__41329),
            .I(port_address_in_2));
    InMux I__10386 (
            .O(N__41326),
            .I(N__41323));
    LocalMux I__10385 (
            .O(N__41323),
            .I(N__41320));
    Odrv4 I__10384 (
            .O(N__41320),
            .I(port_address_in_3));
    InMux I__10383 (
            .O(N__41317),
            .I(N__41314));
    LocalMux I__10382 (
            .O(N__41314),
            .I(port_address_in_6));
    InMux I__10381 (
            .O(N__41311),
            .I(N__41308));
    LocalMux I__10380 (
            .O(N__41308),
            .I(N__41305));
    Span12Mux_v I__10379 (
            .O(N__41305),
            .I(N__41302));
    Odrv12 I__10378 (
            .O(N__41302),
            .I(port_address_in_5));
    CascadeMux I__10377 (
            .O(N__41299),
            .I(N__41296));
    InMux I__10376 (
            .O(N__41296),
            .I(N__41293));
    LocalMux I__10375 (
            .O(N__41293),
            .I(N__41290));
    Span12Mux_s1_h I__10374 (
            .O(N__41290),
            .I(N__41287));
    Odrv12 I__10373 (
            .O(N__41287),
            .I(\this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0 ));
    InMux I__10372 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__10371 (
            .O(N__41281),
            .I(N__41278));
    Span12Mux_s2_h I__10370 (
            .O(N__41278),
            .I(N__41275));
    Span12Mux_v I__10369 (
            .O(N__41275),
            .I(N__41272));
    Odrv12 I__10368 (
            .O(N__41272),
            .I(port_address_in_7));
    InMux I__10367 (
            .O(N__41269),
            .I(N__41266));
    LocalMux I__10366 (
            .O(N__41266),
            .I(N__41263));
    Span4Mux_v I__10365 (
            .O(N__41263),
            .I(N__41260));
    Span4Mux_h I__10364 (
            .O(N__41260),
            .I(N__41256));
    InMux I__10363 (
            .O(N__41259),
            .I(N__41253));
    Sp12to4 I__10362 (
            .O(N__41256),
            .I(N__41248));
    LocalMux I__10361 (
            .O(N__41253),
            .I(N__41248));
    Odrv12 I__10360 (
            .O(N__41248),
            .I(\this_ppu.N_173 ));
    InMux I__10359 (
            .O(N__41245),
            .I(N__41242));
    LocalMux I__10358 (
            .O(N__41242),
            .I(N__41239));
    Span4Mux_v I__10357 (
            .O(N__41239),
            .I(N__41236));
    Odrv4 I__10356 (
            .O(N__41236),
            .I(un1_M_this_ext_address_q_cry_4_THRU_CO));
    IoInMux I__10355 (
            .O(N__41233),
            .I(N__41230));
    LocalMux I__10354 (
            .O(N__41230),
            .I(N__41226));
    InMux I__10353 (
            .O(N__41229),
            .I(N__41223));
    Span4Mux_s2_h I__10352 (
            .O(N__41226),
            .I(N__41219));
    LocalMux I__10351 (
            .O(N__41223),
            .I(N__41216));
    InMux I__10350 (
            .O(N__41222),
            .I(N__41213));
    Span4Mux_h I__10349 (
            .O(N__41219),
            .I(N__41208));
    Span4Mux_h I__10348 (
            .O(N__41216),
            .I(N__41208));
    LocalMux I__10347 (
            .O(N__41213),
            .I(M_this_ext_address_qZ0Z_5));
    Odrv4 I__10346 (
            .O(N__41208),
            .I(M_this_ext_address_qZ0Z_5));
    InMux I__10345 (
            .O(N__41203),
            .I(N__41200));
    LocalMux I__10344 (
            .O(N__41200),
            .I(N__41197));
    Span4Mux_h I__10343 (
            .O(N__41197),
            .I(N__41194));
    Odrv4 I__10342 (
            .O(N__41194),
            .I(un1_M_this_ext_address_q_cry_5_THRU_CO));
    IoInMux I__10341 (
            .O(N__41191),
            .I(N__41188));
    LocalMux I__10340 (
            .O(N__41188),
            .I(N__41185));
    Span4Mux_s2_h I__10339 (
            .O(N__41185),
            .I(N__41181));
    InMux I__10338 (
            .O(N__41184),
            .I(N__41178));
    Span4Mux_v I__10337 (
            .O(N__41181),
            .I(N__41174));
    LocalMux I__10336 (
            .O(N__41178),
            .I(N__41171));
    InMux I__10335 (
            .O(N__41177),
            .I(N__41168));
    Span4Mux_h I__10334 (
            .O(N__41174),
            .I(N__41163));
    Span4Mux_h I__10333 (
            .O(N__41171),
            .I(N__41163));
    LocalMux I__10332 (
            .O(N__41168),
            .I(M_this_ext_address_qZ0Z_6));
    Odrv4 I__10331 (
            .O(N__41163),
            .I(M_this_ext_address_qZ0Z_6));
    InMux I__10330 (
            .O(N__41158),
            .I(N__41155));
    LocalMux I__10329 (
            .O(N__41155),
            .I(N__41152));
    Span4Mux_h I__10328 (
            .O(N__41152),
            .I(N__41149));
    Odrv4 I__10327 (
            .O(N__41149),
            .I(un1_M_this_ext_address_q_cry_6_THRU_CO));
    IoInMux I__10326 (
            .O(N__41146),
            .I(N__41143));
    LocalMux I__10325 (
            .O(N__41143),
            .I(N__41140));
    IoSpan4Mux I__10324 (
            .O(N__41140),
            .I(N__41137));
    Span4Mux_s2_h I__10323 (
            .O(N__41137),
            .I(N__41133));
    CascadeMux I__10322 (
            .O(N__41136),
            .I(N__41130));
    Span4Mux_h I__10321 (
            .O(N__41133),
            .I(N__41127));
    InMux I__10320 (
            .O(N__41130),
            .I(N__41124));
    Sp12to4 I__10319 (
            .O(N__41127),
            .I(N__41121));
    LocalMux I__10318 (
            .O(N__41124),
            .I(N__41117));
    Span12Mux_v I__10317 (
            .O(N__41121),
            .I(N__41114));
    InMux I__10316 (
            .O(N__41120),
            .I(N__41111));
    Span4Mux_h I__10315 (
            .O(N__41117),
            .I(N__41108));
    Odrv12 I__10314 (
            .O(N__41114),
            .I(M_this_ext_address_qZ0Z_7));
    LocalMux I__10313 (
            .O(N__41111),
            .I(M_this_ext_address_qZ0Z_7));
    Odrv4 I__10312 (
            .O(N__41108),
            .I(M_this_ext_address_qZ0Z_7));
    InMux I__10311 (
            .O(N__41101),
            .I(N__41098));
    LocalMux I__10310 (
            .O(N__41098),
            .I(N__41095));
    Odrv4 I__10309 (
            .O(N__41095),
            .I(un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0));
    IoInMux I__10308 (
            .O(N__41092),
            .I(N__41089));
    LocalMux I__10307 (
            .O(N__41089),
            .I(N__41086));
    Span4Mux_s3_v I__10306 (
            .O(N__41086),
            .I(N__41083));
    Span4Mux_h I__10305 (
            .O(N__41083),
            .I(N__41079));
    InMux I__10304 (
            .O(N__41082),
            .I(N__41076));
    Span4Mux_v I__10303 (
            .O(N__41079),
            .I(N__41073));
    LocalMux I__10302 (
            .O(N__41076),
            .I(N__41070));
    Odrv4 I__10301 (
            .O(N__41073),
            .I(M_this_ext_address_qZ0Z_11));
    Odrv12 I__10300 (
            .O(N__41070),
            .I(M_this_ext_address_qZ0Z_11));
    InMux I__10299 (
            .O(N__41065),
            .I(N__41062));
    LocalMux I__10298 (
            .O(N__41062),
            .I(N__41059));
    Odrv4 I__10297 (
            .O(N__41059),
            .I(un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0));
    CascadeMux I__10296 (
            .O(N__41056),
            .I(N__41051));
    InMux I__10295 (
            .O(N__41055),
            .I(N__41048));
    InMux I__10294 (
            .O(N__41054),
            .I(N__41045));
    InMux I__10293 (
            .O(N__41051),
            .I(N__41042));
    LocalMux I__10292 (
            .O(N__41048),
            .I(N__41036));
    LocalMux I__10291 (
            .O(N__41045),
            .I(N__41033));
    LocalMux I__10290 (
            .O(N__41042),
            .I(N__41030));
    InMux I__10289 (
            .O(N__41041),
            .I(N__41026));
    CascadeMux I__10288 (
            .O(N__41040),
            .I(N__41023));
    InMux I__10287 (
            .O(N__41039),
            .I(N__41020));
    Span4Mux_v I__10286 (
            .O(N__41036),
            .I(N__41017));
    Span4Mux_v I__10285 (
            .O(N__41033),
            .I(N__41013));
    Span4Mux_v I__10284 (
            .O(N__41030),
            .I(N__41010));
    InMux I__10283 (
            .O(N__41029),
            .I(N__41007));
    LocalMux I__10282 (
            .O(N__41026),
            .I(N__41004));
    InMux I__10281 (
            .O(N__41023),
            .I(N__41001));
    LocalMux I__10280 (
            .O(N__41020),
            .I(N__40998));
    Span4Mux_v I__10279 (
            .O(N__41017),
            .I(N__40995));
    InMux I__10278 (
            .O(N__41016),
            .I(N__40992));
    Span4Mux_h I__10277 (
            .O(N__41013),
            .I(N__40989));
    Span4Mux_v I__10276 (
            .O(N__41010),
            .I(N__40984));
    LocalMux I__10275 (
            .O(N__41007),
            .I(N__40984));
    Span12Mux_h I__10274 (
            .O(N__41004),
            .I(N__40980));
    LocalMux I__10273 (
            .O(N__41001),
            .I(N__40977));
    Span12Mux_v I__10272 (
            .O(N__40998),
            .I(N__40974));
    Span4Mux_h I__10271 (
            .O(N__40995),
            .I(N__40971));
    LocalMux I__10270 (
            .O(N__40992),
            .I(N__40968));
    Span4Mux_h I__10269 (
            .O(N__40989),
            .I(N__40963));
    Span4Mux_v I__10268 (
            .O(N__40984),
            .I(N__40963));
    InMux I__10267 (
            .O(N__40983),
            .I(N__40960));
    Span12Mux_v I__10266 (
            .O(N__40980),
            .I(N__40957));
    Span12Mux_v I__10265 (
            .O(N__40977),
            .I(N__40954));
    Span12Mux_h I__10264 (
            .O(N__40974),
            .I(N__40943));
    Sp12to4 I__10263 (
            .O(N__40971),
            .I(N__40943));
    Span12Mux_v I__10262 (
            .O(N__40968),
            .I(N__40943));
    Sp12to4 I__10261 (
            .O(N__40963),
            .I(N__40943));
    LocalMux I__10260 (
            .O(N__40960),
            .I(N__40943));
    Odrv12 I__10259 (
            .O(N__40957),
            .I(port_data_c_4));
    Odrv12 I__10258 (
            .O(N__40954),
            .I(port_data_c_4));
    Odrv12 I__10257 (
            .O(N__40943),
            .I(port_data_c_4));
    IoInMux I__10256 (
            .O(N__40936),
            .I(N__40933));
    LocalMux I__10255 (
            .O(N__40933),
            .I(N__40930));
    Span4Mux_s2_h I__10254 (
            .O(N__40930),
            .I(N__40926));
    InMux I__10253 (
            .O(N__40929),
            .I(N__40923));
    Span4Mux_h I__10252 (
            .O(N__40926),
            .I(N__40920));
    LocalMux I__10251 (
            .O(N__40923),
            .I(N__40917));
    Odrv4 I__10250 (
            .O(N__40920),
            .I(M_this_ext_address_qZ0Z_12));
    Odrv12 I__10249 (
            .O(N__40917),
            .I(M_this_ext_address_qZ0Z_12));
    InMux I__10248 (
            .O(N__40912),
            .I(N__40888));
    InMux I__10247 (
            .O(N__40911),
            .I(N__40888));
    InMux I__10246 (
            .O(N__40910),
            .I(N__40888));
    InMux I__10245 (
            .O(N__40909),
            .I(N__40888));
    InMux I__10244 (
            .O(N__40908),
            .I(N__40888));
    InMux I__10243 (
            .O(N__40907),
            .I(N__40888));
    InMux I__10242 (
            .O(N__40906),
            .I(N__40888));
    InMux I__10241 (
            .O(N__40905),
            .I(N__40888));
    LocalMux I__10240 (
            .O(N__40888),
            .I(N__40876));
    InMux I__10239 (
            .O(N__40887),
            .I(N__40869));
    InMux I__10238 (
            .O(N__40886),
            .I(N__40869));
    InMux I__10237 (
            .O(N__40885),
            .I(N__40869));
    InMux I__10236 (
            .O(N__40884),
            .I(N__40856));
    InMux I__10235 (
            .O(N__40883),
            .I(N__40856));
    InMux I__10234 (
            .O(N__40882),
            .I(N__40856));
    InMux I__10233 (
            .O(N__40881),
            .I(N__40856));
    InMux I__10232 (
            .O(N__40880),
            .I(N__40856));
    InMux I__10231 (
            .O(N__40879),
            .I(N__40856));
    Span4Mux_v I__10230 (
            .O(N__40876),
            .I(N__40852));
    LocalMux I__10229 (
            .O(N__40869),
            .I(N__40849));
    LocalMux I__10228 (
            .O(N__40856),
            .I(N__40840));
    InMux I__10227 (
            .O(N__40855),
            .I(N__40837));
    Span4Mux_h I__10226 (
            .O(N__40852),
            .I(N__40831));
    Span4Mux_v I__10225 (
            .O(N__40849),
            .I(N__40831));
    InMux I__10224 (
            .O(N__40848),
            .I(N__40828));
    InMux I__10223 (
            .O(N__40847),
            .I(N__40824));
    InMux I__10222 (
            .O(N__40846),
            .I(N__40821));
    InMux I__10221 (
            .O(N__40845),
            .I(N__40814));
    InMux I__10220 (
            .O(N__40844),
            .I(N__40814));
    InMux I__10219 (
            .O(N__40843),
            .I(N__40811));
    Span4Mux_v I__10218 (
            .O(N__40840),
            .I(N__40806));
    LocalMux I__10217 (
            .O(N__40837),
            .I(N__40806));
    InMux I__10216 (
            .O(N__40836),
            .I(N__40800));
    Span4Mux_v I__10215 (
            .O(N__40831),
            .I(N__40795));
    LocalMux I__10214 (
            .O(N__40828),
            .I(N__40795));
    InMux I__10213 (
            .O(N__40827),
            .I(N__40790));
    LocalMux I__10212 (
            .O(N__40824),
            .I(N__40785));
    LocalMux I__10211 (
            .O(N__40821),
            .I(N__40785));
    InMux I__10210 (
            .O(N__40820),
            .I(N__40782));
    InMux I__10209 (
            .O(N__40819),
            .I(N__40779));
    LocalMux I__10208 (
            .O(N__40814),
            .I(N__40776));
    LocalMux I__10207 (
            .O(N__40811),
            .I(N__40771));
    Span4Mux_h I__10206 (
            .O(N__40806),
            .I(N__40771));
    InMux I__10205 (
            .O(N__40805),
            .I(N__40766));
    InMux I__10204 (
            .O(N__40804),
            .I(N__40766));
    InMux I__10203 (
            .O(N__40803),
            .I(N__40763));
    LocalMux I__10202 (
            .O(N__40800),
            .I(N__40760));
    Span4Mux_h I__10201 (
            .O(N__40795),
            .I(N__40757));
    InMux I__10200 (
            .O(N__40794),
            .I(N__40752));
    InMux I__10199 (
            .O(N__40793),
            .I(N__40752));
    LocalMux I__10198 (
            .O(N__40790),
            .I(N__40739));
    Span4Mux_h I__10197 (
            .O(N__40785),
            .I(N__40739));
    LocalMux I__10196 (
            .O(N__40782),
            .I(N__40739));
    LocalMux I__10195 (
            .O(N__40779),
            .I(N__40739));
    Span4Mux_v I__10194 (
            .O(N__40776),
            .I(N__40739));
    Span4Mux_v I__10193 (
            .O(N__40771),
            .I(N__40739));
    LocalMux I__10192 (
            .O(N__40766),
            .I(N_309_0));
    LocalMux I__10191 (
            .O(N__40763),
            .I(N_309_0));
    Odrv4 I__10190 (
            .O(N__40760),
            .I(N_309_0));
    Odrv4 I__10189 (
            .O(N__40757),
            .I(N_309_0));
    LocalMux I__10188 (
            .O(N__40752),
            .I(N_309_0));
    Odrv4 I__10187 (
            .O(N__40739),
            .I(N_309_0));
    CascadeMux I__10186 (
            .O(N__40726),
            .I(N__40714));
    CascadeMux I__10185 (
            .O(N__40725),
            .I(N__40711));
    CascadeMux I__10184 (
            .O(N__40724),
            .I(N__40707));
    CascadeMux I__10183 (
            .O(N__40723),
            .I(N__40704));
    CascadeMux I__10182 (
            .O(N__40722),
            .I(N__40696));
    CascadeMux I__10181 (
            .O(N__40721),
            .I(N__40693));
    CascadeMux I__10180 (
            .O(N__40720),
            .I(N__40690));
    InMux I__10179 (
            .O(N__40719),
            .I(N__40683));
    InMux I__10178 (
            .O(N__40718),
            .I(N__40683));
    InMux I__10177 (
            .O(N__40717),
            .I(N__40683));
    InMux I__10176 (
            .O(N__40714),
            .I(N__40676));
    InMux I__10175 (
            .O(N__40711),
            .I(N__40676));
    InMux I__10174 (
            .O(N__40710),
            .I(N__40676));
    InMux I__10173 (
            .O(N__40707),
            .I(N__40665));
    InMux I__10172 (
            .O(N__40704),
            .I(N__40665));
    InMux I__10171 (
            .O(N__40703),
            .I(N__40665));
    InMux I__10170 (
            .O(N__40702),
            .I(N__40665));
    InMux I__10169 (
            .O(N__40701),
            .I(N__40665));
    InMux I__10168 (
            .O(N__40700),
            .I(N__40653));
    InMux I__10167 (
            .O(N__40699),
            .I(N__40653));
    InMux I__10166 (
            .O(N__40696),
            .I(N__40653));
    InMux I__10165 (
            .O(N__40693),
            .I(N__40653));
    InMux I__10164 (
            .O(N__40690),
            .I(N__40653));
    LocalMux I__10163 (
            .O(N__40683),
            .I(N__40650));
    LocalMux I__10162 (
            .O(N__40676),
            .I(N__40645));
    LocalMux I__10161 (
            .O(N__40665),
            .I(N__40645));
    CascadeMux I__10160 (
            .O(N__40664),
            .I(N__40642));
    LocalMux I__10159 (
            .O(N__40653),
            .I(N__40639));
    Span4Mux_h I__10158 (
            .O(N__40650),
            .I(N__40636));
    Span4Mux_v I__10157 (
            .O(N__40645),
            .I(N__40633));
    InMux I__10156 (
            .O(N__40642),
            .I(N__40630));
    Span4Mux_v I__10155 (
            .O(N__40639),
            .I(N__40627));
    Span4Mux_v I__10154 (
            .O(N__40636),
            .I(N__40624));
    Span4Mux_h I__10153 (
            .O(N__40633),
            .I(N__40621));
    LocalMux I__10152 (
            .O(N__40630),
            .I(N__40618));
    Odrv4 I__10151 (
            .O(N__40627),
            .I(N_311_0));
    Odrv4 I__10150 (
            .O(N__40624),
            .I(N_311_0));
    Odrv4 I__10149 (
            .O(N__40621),
            .I(N_311_0));
    Odrv4 I__10148 (
            .O(N__40618),
            .I(N_311_0));
    CascadeMux I__10147 (
            .O(N__40609),
            .I(N__40604));
    InMux I__10146 (
            .O(N__40608),
            .I(N__40601));
    InMux I__10145 (
            .O(N__40607),
            .I(N__40595));
    InMux I__10144 (
            .O(N__40604),
            .I(N__40592));
    LocalMux I__10143 (
            .O(N__40601),
            .I(N__40589));
    InMux I__10142 (
            .O(N__40600),
            .I(N__40586));
    InMux I__10141 (
            .O(N__40599),
            .I(N__40583));
    InMux I__10140 (
            .O(N__40598),
            .I(N__40579));
    LocalMux I__10139 (
            .O(N__40595),
            .I(N__40576));
    LocalMux I__10138 (
            .O(N__40592),
            .I(N__40571));
    Span4Mux_h I__10137 (
            .O(N__40589),
            .I(N__40566));
    LocalMux I__10136 (
            .O(N__40586),
            .I(N__40566));
    LocalMux I__10135 (
            .O(N__40583),
            .I(N__40563));
    CascadeMux I__10134 (
            .O(N__40582),
            .I(N__40560));
    LocalMux I__10133 (
            .O(N__40579),
            .I(N__40557));
    Span4Mux_h I__10132 (
            .O(N__40576),
            .I(N__40554));
    InMux I__10131 (
            .O(N__40575),
            .I(N__40551));
    InMux I__10130 (
            .O(N__40574),
            .I(N__40548));
    Span4Mux_v I__10129 (
            .O(N__40571),
            .I(N__40545));
    Span4Mux_v I__10128 (
            .O(N__40566),
            .I(N__40540));
    Span4Mux_v I__10127 (
            .O(N__40563),
            .I(N__40540));
    InMux I__10126 (
            .O(N__40560),
            .I(N__40537));
    Span12Mux_v I__10125 (
            .O(N__40557),
            .I(N__40534));
    Sp12to4 I__10124 (
            .O(N__40554),
            .I(N__40527));
    LocalMux I__10123 (
            .O(N__40551),
            .I(N__40527));
    LocalMux I__10122 (
            .O(N__40548),
            .I(N__40527));
    Sp12to4 I__10121 (
            .O(N__40545),
            .I(N__40522));
    Sp12to4 I__10120 (
            .O(N__40540),
            .I(N__40522));
    LocalMux I__10119 (
            .O(N__40537),
            .I(N__40519));
    Span12Mux_h I__10118 (
            .O(N__40534),
            .I(N__40516));
    Span12Mux_v I__10117 (
            .O(N__40527),
            .I(N__40513));
    Span12Mux_h I__10116 (
            .O(N__40522),
            .I(N__40508));
    Span12Mux_v I__10115 (
            .O(N__40519),
            .I(N__40508));
    Odrv12 I__10114 (
            .O(N__40516),
            .I(port_data_c_5));
    Odrv12 I__10113 (
            .O(N__40513),
            .I(port_data_c_5));
    Odrv12 I__10112 (
            .O(N__40508),
            .I(port_data_c_5));
    InMux I__10111 (
            .O(N__40501),
            .I(N__40498));
    LocalMux I__10110 (
            .O(N__40498),
            .I(N__40495));
    Odrv4 I__10109 (
            .O(N__40495),
            .I(un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0));
    IoInMux I__10108 (
            .O(N__40492),
            .I(N__40489));
    LocalMux I__10107 (
            .O(N__40489),
            .I(N__40485));
    CascadeMux I__10106 (
            .O(N__40488),
            .I(N__40482));
    IoSpan4Mux I__10105 (
            .O(N__40485),
            .I(N__40479));
    InMux I__10104 (
            .O(N__40482),
            .I(N__40476));
    Span4Mux_s3_h I__10103 (
            .O(N__40479),
            .I(N__40473));
    LocalMux I__10102 (
            .O(N__40476),
            .I(N__40470));
    Odrv4 I__10101 (
            .O(N__40473),
            .I(M_this_ext_address_qZ0Z_13));
    Odrv4 I__10100 (
            .O(N__40470),
            .I(M_this_ext_address_qZ0Z_13));
    ClkMux I__10099 (
            .O(N__40465),
            .I(N__39928));
    ClkMux I__10098 (
            .O(N__40464),
            .I(N__39928));
    ClkMux I__10097 (
            .O(N__40463),
            .I(N__39928));
    ClkMux I__10096 (
            .O(N__40462),
            .I(N__39928));
    ClkMux I__10095 (
            .O(N__40461),
            .I(N__39928));
    ClkMux I__10094 (
            .O(N__40460),
            .I(N__39928));
    ClkMux I__10093 (
            .O(N__40459),
            .I(N__39928));
    ClkMux I__10092 (
            .O(N__40458),
            .I(N__39928));
    ClkMux I__10091 (
            .O(N__40457),
            .I(N__39928));
    ClkMux I__10090 (
            .O(N__40456),
            .I(N__39928));
    ClkMux I__10089 (
            .O(N__40455),
            .I(N__39928));
    ClkMux I__10088 (
            .O(N__40454),
            .I(N__39928));
    ClkMux I__10087 (
            .O(N__40453),
            .I(N__39928));
    ClkMux I__10086 (
            .O(N__40452),
            .I(N__39928));
    ClkMux I__10085 (
            .O(N__40451),
            .I(N__39928));
    ClkMux I__10084 (
            .O(N__40450),
            .I(N__39928));
    ClkMux I__10083 (
            .O(N__40449),
            .I(N__39928));
    ClkMux I__10082 (
            .O(N__40448),
            .I(N__39928));
    ClkMux I__10081 (
            .O(N__40447),
            .I(N__39928));
    ClkMux I__10080 (
            .O(N__40446),
            .I(N__39928));
    ClkMux I__10079 (
            .O(N__40445),
            .I(N__39928));
    ClkMux I__10078 (
            .O(N__40444),
            .I(N__39928));
    ClkMux I__10077 (
            .O(N__40443),
            .I(N__39928));
    ClkMux I__10076 (
            .O(N__40442),
            .I(N__39928));
    ClkMux I__10075 (
            .O(N__40441),
            .I(N__39928));
    ClkMux I__10074 (
            .O(N__40440),
            .I(N__39928));
    ClkMux I__10073 (
            .O(N__40439),
            .I(N__39928));
    ClkMux I__10072 (
            .O(N__40438),
            .I(N__39928));
    ClkMux I__10071 (
            .O(N__40437),
            .I(N__39928));
    ClkMux I__10070 (
            .O(N__40436),
            .I(N__39928));
    ClkMux I__10069 (
            .O(N__40435),
            .I(N__39928));
    ClkMux I__10068 (
            .O(N__40434),
            .I(N__39928));
    ClkMux I__10067 (
            .O(N__40433),
            .I(N__39928));
    ClkMux I__10066 (
            .O(N__40432),
            .I(N__39928));
    ClkMux I__10065 (
            .O(N__40431),
            .I(N__39928));
    ClkMux I__10064 (
            .O(N__40430),
            .I(N__39928));
    ClkMux I__10063 (
            .O(N__40429),
            .I(N__39928));
    ClkMux I__10062 (
            .O(N__40428),
            .I(N__39928));
    ClkMux I__10061 (
            .O(N__40427),
            .I(N__39928));
    ClkMux I__10060 (
            .O(N__40426),
            .I(N__39928));
    ClkMux I__10059 (
            .O(N__40425),
            .I(N__39928));
    ClkMux I__10058 (
            .O(N__40424),
            .I(N__39928));
    ClkMux I__10057 (
            .O(N__40423),
            .I(N__39928));
    ClkMux I__10056 (
            .O(N__40422),
            .I(N__39928));
    ClkMux I__10055 (
            .O(N__40421),
            .I(N__39928));
    ClkMux I__10054 (
            .O(N__40420),
            .I(N__39928));
    ClkMux I__10053 (
            .O(N__40419),
            .I(N__39928));
    ClkMux I__10052 (
            .O(N__40418),
            .I(N__39928));
    ClkMux I__10051 (
            .O(N__40417),
            .I(N__39928));
    ClkMux I__10050 (
            .O(N__40416),
            .I(N__39928));
    ClkMux I__10049 (
            .O(N__40415),
            .I(N__39928));
    ClkMux I__10048 (
            .O(N__40414),
            .I(N__39928));
    ClkMux I__10047 (
            .O(N__40413),
            .I(N__39928));
    ClkMux I__10046 (
            .O(N__40412),
            .I(N__39928));
    ClkMux I__10045 (
            .O(N__40411),
            .I(N__39928));
    ClkMux I__10044 (
            .O(N__40410),
            .I(N__39928));
    ClkMux I__10043 (
            .O(N__40409),
            .I(N__39928));
    ClkMux I__10042 (
            .O(N__40408),
            .I(N__39928));
    ClkMux I__10041 (
            .O(N__40407),
            .I(N__39928));
    ClkMux I__10040 (
            .O(N__40406),
            .I(N__39928));
    ClkMux I__10039 (
            .O(N__40405),
            .I(N__39928));
    ClkMux I__10038 (
            .O(N__40404),
            .I(N__39928));
    ClkMux I__10037 (
            .O(N__40403),
            .I(N__39928));
    ClkMux I__10036 (
            .O(N__40402),
            .I(N__39928));
    ClkMux I__10035 (
            .O(N__40401),
            .I(N__39928));
    ClkMux I__10034 (
            .O(N__40400),
            .I(N__39928));
    ClkMux I__10033 (
            .O(N__40399),
            .I(N__39928));
    ClkMux I__10032 (
            .O(N__40398),
            .I(N__39928));
    ClkMux I__10031 (
            .O(N__40397),
            .I(N__39928));
    ClkMux I__10030 (
            .O(N__40396),
            .I(N__39928));
    ClkMux I__10029 (
            .O(N__40395),
            .I(N__39928));
    ClkMux I__10028 (
            .O(N__40394),
            .I(N__39928));
    ClkMux I__10027 (
            .O(N__40393),
            .I(N__39928));
    ClkMux I__10026 (
            .O(N__40392),
            .I(N__39928));
    ClkMux I__10025 (
            .O(N__40391),
            .I(N__39928));
    ClkMux I__10024 (
            .O(N__40390),
            .I(N__39928));
    ClkMux I__10023 (
            .O(N__40389),
            .I(N__39928));
    ClkMux I__10022 (
            .O(N__40388),
            .I(N__39928));
    ClkMux I__10021 (
            .O(N__40387),
            .I(N__39928));
    ClkMux I__10020 (
            .O(N__40386),
            .I(N__39928));
    ClkMux I__10019 (
            .O(N__40385),
            .I(N__39928));
    ClkMux I__10018 (
            .O(N__40384),
            .I(N__39928));
    ClkMux I__10017 (
            .O(N__40383),
            .I(N__39928));
    ClkMux I__10016 (
            .O(N__40382),
            .I(N__39928));
    ClkMux I__10015 (
            .O(N__40381),
            .I(N__39928));
    ClkMux I__10014 (
            .O(N__40380),
            .I(N__39928));
    ClkMux I__10013 (
            .O(N__40379),
            .I(N__39928));
    ClkMux I__10012 (
            .O(N__40378),
            .I(N__39928));
    ClkMux I__10011 (
            .O(N__40377),
            .I(N__39928));
    ClkMux I__10010 (
            .O(N__40376),
            .I(N__39928));
    ClkMux I__10009 (
            .O(N__40375),
            .I(N__39928));
    ClkMux I__10008 (
            .O(N__40374),
            .I(N__39928));
    ClkMux I__10007 (
            .O(N__40373),
            .I(N__39928));
    ClkMux I__10006 (
            .O(N__40372),
            .I(N__39928));
    ClkMux I__10005 (
            .O(N__40371),
            .I(N__39928));
    ClkMux I__10004 (
            .O(N__40370),
            .I(N__39928));
    ClkMux I__10003 (
            .O(N__40369),
            .I(N__39928));
    ClkMux I__10002 (
            .O(N__40368),
            .I(N__39928));
    ClkMux I__10001 (
            .O(N__40367),
            .I(N__39928));
    ClkMux I__10000 (
            .O(N__40366),
            .I(N__39928));
    ClkMux I__9999 (
            .O(N__40365),
            .I(N__39928));
    ClkMux I__9998 (
            .O(N__40364),
            .I(N__39928));
    ClkMux I__9997 (
            .O(N__40363),
            .I(N__39928));
    ClkMux I__9996 (
            .O(N__40362),
            .I(N__39928));
    ClkMux I__9995 (
            .O(N__40361),
            .I(N__39928));
    ClkMux I__9994 (
            .O(N__40360),
            .I(N__39928));
    ClkMux I__9993 (
            .O(N__40359),
            .I(N__39928));
    ClkMux I__9992 (
            .O(N__40358),
            .I(N__39928));
    ClkMux I__9991 (
            .O(N__40357),
            .I(N__39928));
    ClkMux I__9990 (
            .O(N__40356),
            .I(N__39928));
    ClkMux I__9989 (
            .O(N__40355),
            .I(N__39928));
    ClkMux I__9988 (
            .O(N__40354),
            .I(N__39928));
    ClkMux I__9987 (
            .O(N__40353),
            .I(N__39928));
    ClkMux I__9986 (
            .O(N__40352),
            .I(N__39928));
    ClkMux I__9985 (
            .O(N__40351),
            .I(N__39928));
    ClkMux I__9984 (
            .O(N__40350),
            .I(N__39928));
    ClkMux I__9983 (
            .O(N__40349),
            .I(N__39928));
    ClkMux I__9982 (
            .O(N__40348),
            .I(N__39928));
    ClkMux I__9981 (
            .O(N__40347),
            .I(N__39928));
    ClkMux I__9980 (
            .O(N__40346),
            .I(N__39928));
    ClkMux I__9979 (
            .O(N__40345),
            .I(N__39928));
    ClkMux I__9978 (
            .O(N__40344),
            .I(N__39928));
    ClkMux I__9977 (
            .O(N__40343),
            .I(N__39928));
    ClkMux I__9976 (
            .O(N__40342),
            .I(N__39928));
    ClkMux I__9975 (
            .O(N__40341),
            .I(N__39928));
    ClkMux I__9974 (
            .O(N__40340),
            .I(N__39928));
    ClkMux I__9973 (
            .O(N__40339),
            .I(N__39928));
    ClkMux I__9972 (
            .O(N__40338),
            .I(N__39928));
    ClkMux I__9971 (
            .O(N__40337),
            .I(N__39928));
    ClkMux I__9970 (
            .O(N__40336),
            .I(N__39928));
    ClkMux I__9969 (
            .O(N__40335),
            .I(N__39928));
    ClkMux I__9968 (
            .O(N__40334),
            .I(N__39928));
    ClkMux I__9967 (
            .O(N__40333),
            .I(N__39928));
    ClkMux I__9966 (
            .O(N__40332),
            .I(N__39928));
    ClkMux I__9965 (
            .O(N__40331),
            .I(N__39928));
    ClkMux I__9964 (
            .O(N__40330),
            .I(N__39928));
    ClkMux I__9963 (
            .O(N__40329),
            .I(N__39928));
    ClkMux I__9962 (
            .O(N__40328),
            .I(N__39928));
    ClkMux I__9961 (
            .O(N__40327),
            .I(N__39928));
    ClkMux I__9960 (
            .O(N__40326),
            .I(N__39928));
    ClkMux I__9959 (
            .O(N__40325),
            .I(N__39928));
    ClkMux I__9958 (
            .O(N__40324),
            .I(N__39928));
    ClkMux I__9957 (
            .O(N__40323),
            .I(N__39928));
    ClkMux I__9956 (
            .O(N__40322),
            .I(N__39928));
    ClkMux I__9955 (
            .O(N__40321),
            .I(N__39928));
    ClkMux I__9954 (
            .O(N__40320),
            .I(N__39928));
    ClkMux I__9953 (
            .O(N__40319),
            .I(N__39928));
    ClkMux I__9952 (
            .O(N__40318),
            .I(N__39928));
    ClkMux I__9951 (
            .O(N__40317),
            .I(N__39928));
    ClkMux I__9950 (
            .O(N__40316),
            .I(N__39928));
    ClkMux I__9949 (
            .O(N__40315),
            .I(N__39928));
    ClkMux I__9948 (
            .O(N__40314),
            .I(N__39928));
    ClkMux I__9947 (
            .O(N__40313),
            .I(N__39928));
    ClkMux I__9946 (
            .O(N__40312),
            .I(N__39928));
    ClkMux I__9945 (
            .O(N__40311),
            .I(N__39928));
    ClkMux I__9944 (
            .O(N__40310),
            .I(N__39928));
    ClkMux I__9943 (
            .O(N__40309),
            .I(N__39928));
    ClkMux I__9942 (
            .O(N__40308),
            .I(N__39928));
    ClkMux I__9941 (
            .O(N__40307),
            .I(N__39928));
    ClkMux I__9940 (
            .O(N__40306),
            .I(N__39928));
    ClkMux I__9939 (
            .O(N__40305),
            .I(N__39928));
    ClkMux I__9938 (
            .O(N__40304),
            .I(N__39928));
    ClkMux I__9937 (
            .O(N__40303),
            .I(N__39928));
    ClkMux I__9936 (
            .O(N__40302),
            .I(N__39928));
    ClkMux I__9935 (
            .O(N__40301),
            .I(N__39928));
    ClkMux I__9934 (
            .O(N__40300),
            .I(N__39928));
    ClkMux I__9933 (
            .O(N__40299),
            .I(N__39928));
    ClkMux I__9932 (
            .O(N__40298),
            .I(N__39928));
    ClkMux I__9931 (
            .O(N__40297),
            .I(N__39928));
    ClkMux I__9930 (
            .O(N__40296),
            .I(N__39928));
    ClkMux I__9929 (
            .O(N__40295),
            .I(N__39928));
    ClkMux I__9928 (
            .O(N__40294),
            .I(N__39928));
    ClkMux I__9927 (
            .O(N__40293),
            .I(N__39928));
    ClkMux I__9926 (
            .O(N__40292),
            .I(N__39928));
    ClkMux I__9925 (
            .O(N__40291),
            .I(N__39928));
    ClkMux I__9924 (
            .O(N__40290),
            .I(N__39928));
    ClkMux I__9923 (
            .O(N__40289),
            .I(N__39928));
    ClkMux I__9922 (
            .O(N__40288),
            .I(N__39928));
    ClkMux I__9921 (
            .O(N__40287),
            .I(N__39928));
    GlobalMux I__9920 (
            .O(N__39928),
            .I(N__39925));
    gio2CtrlBuf I__9919 (
            .O(N__39925),
            .I(clk_0_c_g));
    CascadeMux I__9918 (
            .O(N__39922),
            .I(N__39916));
    CascadeMux I__9917 (
            .O(N__39921),
            .I(N__39905));
    CascadeMux I__9916 (
            .O(N__39920),
            .I(N__39898));
    CascadeMux I__9915 (
            .O(N__39919),
            .I(N__39886));
    InMux I__9914 (
            .O(N__39916),
            .I(N__39878));
    InMux I__9913 (
            .O(N__39915),
            .I(N__39875));
    InMux I__9912 (
            .O(N__39914),
            .I(N__39872));
    InMux I__9911 (
            .O(N__39913),
            .I(N__39869));
    InMux I__9910 (
            .O(N__39912),
            .I(N__39866));
    InMux I__9909 (
            .O(N__39911),
            .I(N__39863));
    InMux I__9908 (
            .O(N__39910),
            .I(N__39858));
    InMux I__9907 (
            .O(N__39909),
            .I(N__39858));
    InMux I__9906 (
            .O(N__39908),
            .I(N__39855));
    InMux I__9905 (
            .O(N__39905),
            .I(N__39852));
    InMux I__9904 (
            .O(N__39904),
            .I(N__39849));
    InMux I__9903 (
            .O(N__39903),
            .I(N__39846));
    InMux I__9902 (
            .O(N__39902),
            .I(N__39841));
    InMux I__9901 (
            .O(N__39901),
            .I(N__39841));
    InMux I__9900 (
            .O(N__39898),
            .I(N__39838));
    InMux I__9899 (
            .O(N__39897),
            .I(N__39835));
    InMux I__9898 (
            .O(N__39896),
            .I(N__39832));
    InMux I__9897 (
            .O(N__39895),
            .I(N__39829));
    InMux I__9896 (
            .O(N__39894),
            .I(N__39826));
    InMux I__9895 (
            .O(N__39893),
            .I(N__39821));
    InMux I__9894 (
            .O(N__39892),
            .I(N__39821));
    InMux I__9893 (
            .O(N__39891),
            .I(N__39818));
    InMux I__9892 (
            .O(N__39890),
            .I(N__39815));
    InMux I__9891 (
            .O(N__39889),
            .I(N__39812));
    InMux I__9890 (
            .O(N__39886),
            .I(N__39809));
    InMux I__9889 (
            .O(N__39885),
            .I(N__39804));
    InMux I__9888 (
            .O(N__39884),
            .I(N__39804));
    InMux I__9887 (
            .O(N__39883),
            .I(N__39801));
    InMux I__9886 (
            .O(N__39882),
            .I(N__39796));
    InMux I__9885 (
            .O(N__39881),
            .I(N__39796));
    LocalMux I__9884 (
            .O(N__39878),
            .I(N__39751));
    LocalMux I__9883 (
            .O(N__39875),
            .I(N__39748));
    LocalMux I__9882 (
            .O(N__39872),
            .I(N__39745));
    LocalMux I__9881 (
            .O(N__39869),
            .I(N__39742));
    LocalMux I__9880 (
            .O(N__39866),
            .I(N__39739));
    LocalMux I__9879 (
            .O(N__39863),
            .I(N__39736));
    LocalMux I__9878 (
            .O(N__39858),
            .I(N__39733));
    LocalMux I__9877 (
            .O(N__39855),
            .I(N__39730));
    LocalMux I__9876 (
            .O(N__39852),
            .I(N__39727));
    LocalMux I__9875 (
            .O(N__39849),
            .I(N__39724));
    LocalMux I__9874 (
            .O(N__39846),
            .I(N__39721));
    LocalMux I__9873 (
            .O(N__39841),
            .I(N__39718));
    LocalMux I__9872 (
            .O(N__39838),
            .I(N__39715));
    LocalMux I__9871 (
            .O(N__39835),
            .I(N__39712));
    LocalMux I__9870 (
            .O(N__39832),
            .I(N__39709));
    LocalMux I__9869 (
            .O(N__39829),
            .I(N__39706));
    LocalMux I__9868 (
            .O(N__39826),
            .I(N__39703));
    LocalMux I__9867 (
            .O(N__39821),
            .I(N__39700));
    LocalMux I__9866 (
            .O(N__39818),
            .I(N__39697));
    LocalMux I__9865 (
            .O(N__39815),
            .I(N__39694));
    LocalMux I__9864 (
            .O(N__39812),
            .I(N__39691));
    LocalMux I__9863 (
            .O(N__39809),
            .I(N__39688));
    LocalMux I__9862 (
            .O(N__39804),
            .I(N__39685));
    LocalMux I__9861 (
            .O(N__39801),
            .I(N__39682));
    LocalMux I__9860 (
            .O(N__39796),
            .I(N__39679));
    SRMux I__9859 (
            .O(N__39795),
            .I(N__39544));
    SRMux I__9858 (
            .O(N__39794),
            .I(N__39544));
    SRMux I__9857 (
            .O(N__39793),
            .I(N__39544));
    SRMux I__9856 (
            .O(N__39792),
            .I(N__39544));
    SRMux I__9855 (
            .O(N__39791),
            .I(N__39544));
    SRMux I__9854 (
            .O(N__39790),
            .I(N__39544));
    SRMux I__9853 (
            .O(N__39789),
            .I(N__39544));
    SRMux I__9852 (
            .O(N__39788),
            .I(N__39544));
    SRMux I__9851 (
            .O(N__39787),
            .I(N__39544));
    SRMux I__9850 (
            .O(N__39786),
            .I(N__39544));
    SRMux I__9849 (
            .O(N__39785),
            .I(N__39544));
    SRMux I__9848 (
            .O(N__39784),
            .I(N__39544));
    SRMux I__9847 (
            .O(N__39783),
            .I(N__39544));
    SRMux I__9846 (
            .O(N__39782),
            .I(N__39544));
    SRMux I__9845 (
            .O(N__39781),
            .I(N__39544));
    SRMux I__9844 (
            .O(N__39780),
            .I(N__39544));
    SRMux I__9843 (
            .O(N__39779),
            .I(N__39544));
    SRMux I__9842 (
            .O(N__39778),
            .I(N__39544));
    SRMux I__9841 (
            .O(N__39777),
            .I(N__39544));
    SRMux I__9840 (
            .O(N__39776),
            .I(N__39544));
    SRMux I__9839 (
            .O(N__39775),
            .I(N__39544));
    SRMux I__9838 (
            .O(N__39774),
            .I(N__39544));
    SRMux I__9837 (
            .O(N__39773),
            .I(N__39544));
    SRMux I__9836 (
            .O(N__39772),
            .I(N__39544));
    SRMux I__9835 (
            .O(N__39771),
            .I(N__39544));
    SRMux I__9834 (
            .O(N__39770),
            .I(N__39544));
    SRMux I__9833 (
            .O(N__39769),
            .I(N__39544));
    SRMux I__9832 (
            .O(N__39768),
            .I(N__39544));
    SRMux I__9831 (
            .O(N__39767),
            .I(N__39544));
    SRMux I__9830 (
            .O(N__39766),
            .I(N__39544));
    SRMux I__9829 (
            .O(N__39765),
            .I(N__39544));
    SRMux I__9828 (
            .O(N__39764),
            .I(N__39544));
    SRMux I__9827 (
            .O(N__39763),
            .I(N__39544));
    SRMux I__9826 (
            .O(N__39762),
            .I(N__39544));
    SRMux I__9825 (
            .O(N__39761),
            .I(N__39544));
    SRMux I__9824 (
            .O(N__39760),
            .I(N__39544));
    SRMux I__9823 (
            .O(N__39759),
            .I(N__39544));
    SRMux I__9822 (
            .O(N__39758),
            .I(N__39544));
    SRMux I__9821 (
            .O(N__39757),
            .I(N__39544));
    SRMux I__9820 (
            .O(N__39756),
            .I(N__39544));
    SRMux I__9819 (
            .O(N__39755),
            .I(N__39544));
    SRMux I__9818 (
            .O(N__39754),
            .I(N__39544));
    Glb2LocalMux I__9817 (
            .O(N__39751),
            .I(N__39544));
    Glb2LocalMux I__9816 (
            .O(N__39748),
            .I(N__39544));
    Glb2LocalMux I__9815 (
            .O(N__39745),
            .I(N__39544));
    Glb2LocalMux I__9814 (
            .O(N__39742),
            .I(N__39544));
    Glb2LocalMux I__9813 (
            .O(N__39739),
            .I(N__39544));
    Glb2LocalMux I__9812 (
            .O(N__39736),
            .I(N__39544));
    Glb2LocalMux I__9811 (
            .O(N__39733),
            .I(N__39544));
    Glb2LocalMux I__9810 (
            .O(N__39730),
            .I(N__39544));
    Glb2LocalMux I__9809 (
            .O(N__39727),
            .I(N__39544));
    Glb2LocalMux I__9808 (
            .O(N__39724),
            .I(N__39544));
    Glb2LocalMux I__9807 (
            .O(N__39721),
            .I(N__39544));
    Glb2LocalMux I__9806 (
            .O(N__39718),
            .I(N__39544));
    Glb2LocalMux I__9805 (
            .O(N__39715),
            .I(N__39544));
    Glb2LocalMux I__9804 (
            .O(N__39712),
            .I(N__39544));
    Glb2LocalMux I__9803 (
            .O(N__39709),
            .I(N__39544));
    Glb2LocalMux I__9802 (
            .O(N__39706),
            .I(N__39544));
    Glb2LocalMux I__9801 (
            .O(N__39703),
            .I(N__39544));
    Glb2LocalMux I__9800 (
            .O(N__39700),
            .I(N__39544));
    Glb2LocalMux I__9799 (
            .O(N__39697),
            .I(N__39544));
    Glb2LocalMux I__9798 (
            .O(N__39694),
            .I(N__39544));
    Glb2LocalMux I__9797 (
            .O(N__39691),
            .I(N__39544));
    Glb2LocalMux I__9796 (
            .O(N__39688),
            .I(N__39544));
    Glb2LocalMux I__9795 (
            .O(N__39685),
            .I(N__39544));
    Glb2LocalMux I__9794 (
            .O(N__39682),
            .I(N__39544));
    Glb2LocalMux I__9793 (
            .O(N__39679),
            .I(N__39544));
    GlobalMux I__9792 (
            .O(N__39544),
            .I(N__39541));
    gio2CtrlBuf I__9791 (
            .O(N__39541),
            .I(M_this_reset_cond_out_g_0));
    InMux I__9790 (
            .O(N__39538),
            .I(N__39535));
    LocalMux I__9789 (
            .O(N__39535),
            .I(N__39532));
    Odrv4 I__9788 (
            .O(N__39532),
            .I(M_this_oam_ram_read_data_12));
    InMux I__9787 (
            .O(N__39529),
            .I(N__39526));
    LocalMux I__9786 (
            .O(N__39526),
            .I(N__39523));
    Span4Mux_v I__9785 (
            .O(N__39523),
            .I(N__39520));
    Odrv4 I__9784 (
            .O(N__39520),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_12 ));
    InMux I__9783 (
            .O(N__39517),
            .I(N__39513));
    CascadeMux I__9782 (
            .O(N__39516),
            .I(N__39510));
    LocalMux I__9781 (
            .O(N__39513),
            .I(N__39507));
    InMux I__9780 (
            .O(N__39510),
            .I(N__39502));
    Span4Mux_h I__9779 (
            .O(N__39507),
            .I(N__39499));
    InMux I__9778 (
            .O(N__39506),
            .I(N__39494));
    CascadeMux I__9777 (
            .O(N__39505),
            .I(N__39491));
    LocalMux I__9776 (
            .O(N__39502),
            .I(N__39488));
    Span4Mux_v I__9775 (
            .O(N__39499),
            .I(N__39485));
    InMux I__9774 (
            .O(N__39498),
            .I(N__39482));
    InMux I__9773 (
            .O(N__39497),
            .I(N__39479));
    LocalMux I__9772 (
            .O(N__39494),
            .I(N__39475));
    InMux I__9771 (
            .O(N__39491),
            .I(N__39472));
    Span4Mux_v I__9770 (
            .O(N__39488),
            .I(N__39469));
    Span4Mux_h I__9769 (
            .O(N__39485),
            .I(N__39464));
    LocalMux I__9768 (
            .O(N__39482),
            .I(N__39464));
    LocalMux I__9767 (
            .O(N__39479),
            .I(N__39461));
    InMux I__9766 (
            .O(N__39478),
            .I(N__39458));
    Span4Mux_v I__9765 (
            .O(N__39475),
            .I(N__39455));
    LocalMux I__9764 (
            .O(N__39472),
            .I(N__39451));
    Span4Mux_v I__9763 (
            .O(N__39469),
            .I(N__39448));
    Span4Mux_h I__9762 (
            .O(N__39464),
            .I(N__39441));
    Span4Mux_v I__9761 (
            .O(N__39461),
            .I(N__39441));
    LocalMux I__9760 (
            .O(N__39458),
            .I(N__39441));
    Sp12to4 I__9759 (
            .O(N__39455),
            .I(N__39437));
    InMux I__9758 (
            .O(N__39454),
            .I(N__39434));
    Span4Mux_h I__9757 (
            .O(N__39451),
            .I(N__39431));
    Span4Mux_v I__9756 (
            .O(N__39448),
            .I(N__39426));
    Span4Mux_h I__9755 (
            .O(N__39441),
            .I(N__39426));
    InMux I__9754 (
            .O(N__39440),
            .I(N__39423));
    Span12Mux_h I__9753 (
            .O(N__39437),
            .I(N__39420));
    LocalMux I__9752 (
            .O(N__39434),
            .I(N__39417));
    Span4Mux_v I__9751 (
            .O(N__39431),
            .I(N__39414));
    Span4Mux_h I__9750 (
            .O(N__39426),
            .I(N__39411));
    LocalMux I__9749 (
            .O(N__39423),
            .I(N__39408));
    Span12Mux_v I__9748 (
            .O(N__39420),
            .I(N__39405));
    Span12Mux_h I__9747 (
            .O(N__39417),
            .I(N__39402));
    Span4Mux_v I__9746 (
            .O(N__39414),
            .I(N__39399));
    Span4Mux_v I__9745 (
            .O(N__39411),
            .I(N__39394));
    Span4Mux_h I__9744 (
            .O(N__39408),
            .I(N__39394));
    Odrv12 I__9743 (
            .O(N__39405),
            .I(port_data_c_3));
    Odrv12 I__9742 (
            .O(N__39402),
            .I(port_data_c_3));
    Odrv4 I__9741 (
            .O(N__39399),
            .I(port_data_c_3));
    Odrv4 I__9740 (
            .O(N__39394),
            .I(port_data_c_3));
    CEMux I__9739 (
            .O(N__39385),
            .I(N__39381));
    CEMux I__9738 (
            .O(N__39384),
            .I(N__39378));
    LocalMux I__9737 (
            .O(N__39381),
            .I(N__39365));
    LocalMux I__9736 (
            .O(N__39378),
            .I(N__39362));
    InMux I__9735 (
            .O(N__39377),
            .I(N__39355));
    InMux I__9734 (
            .O(N__39376),
            .I(N__39355));
    InMux I__9733 (
            .O(N__39375),
            .I(N__39355));
    InMux I__9732 (
            .O(N__39374),
            .I(N__39350));
    InMux I__9731 (
            .O(N__39373),
            .I(N__39350));
    InMux I__9730 (
            .O(N__39372),
            .I(N__39343));
    InMux I__9729 (
            .O(N__39371),
            .I(N__39336));
    InMux I__9728 (
            .O(N__39370),
            .I(N__39336));
    InMux I__9727 (
            .O(N__39369),
            .I(N__39336));
    InMux I__9726 (
            .O(N__39368),
            .I(N__39330));
    Span4Mux_h I__9725 (
            .O(N__39365),
            .I(N__39325));
    Span4Mux_v I__9724 (
            .O(N__39362),
            .I(N__39320));
    LocalMux I__9723 (
            .O(N__39355),
            .I(N__39320));
    LocalMux I__9722 (
            .O(N__39350),
            .I(N__39309));
    InMux I__9721 (
            .O(N__39349),
            .I(N__39298));
    InMux I__9720 (
            .O(N__39348),
            .I(N__39298));
    InMux I__9719 (
            .O(N__39347),
            .I(N__39298));
    InMux I__9718 (
            .O(N__39346),
            .I(N__39298));
    LocalMux I__9717 (
            .O(N__39343),
            .I(N__39293));
    LocalMux I__9716 (
            .O(N__39336),
            .I(N__39293));
    InMux I__9715 (
            .O(N__39335),
            .I(N__39286));
    InMux I__9714 (
            .O(N__39334),
            .I(N__39286));
    InMux I__9713 (
            .O(N__39333),
            .I(N__39286));
    LocalMux I__9712 (
            .O(N__39330),
            .I(N__39283));
    InMux I__9711 (
            .O(N__39329),
            .I(N__39280));
    InMux I__9710 (
            .O(N__39328),
            .I(N__39277));
    Span4Mux_v I__9709 (
            .O(N__39325),
            .I(N__39272));
    Span4Mux_h I__9708 (
            .O(N__39320),
            .I(N__39272));
    InMux I__9707 (
            .O(N__39319),
            .I(N__39266));
    InMux I__9706 (
            .O(N__39318),
            .I(N__39263));
    InMux I__9705 (
            .O(N__39317),
            .I(N__39258));
    InMux I__9704 (
            .O(N__39316),
            .I(N__39258));
    InMux I__9703 (
            .O(N__39315),
            .I(N__39255));
    InMux I__9702 (
            .O(N__39314),
            .I(N__39252));
    InMux I__9701 (
            .O(N__39313),
            .I(N__39247));
    InMux I__9700 (
            .O(N__39312),
            .I(N__39247));
    Span4Mux_h I__9699 (
            .O(N__39309),
            .I(N__39244));
    InMux I__9698 (
            .O(N__39308),
            .I(N__39241));
    InMux I__9697 (
            .O(N__39307),
            .I(N__39238));
    LocalMux I__9696 (
            .O(N__39298),
            .I(N__39231));
    Span4Mux_v I__9695 (
            .O(N__39293),
            .I(N__39231));
    LocalMux I__9694 (
            .O(N__39286),
            .I(N__39231));
    Span4Mux_v I__9693 (
            .O(N__39283),
            .I(N__39224));
    LocalMux I__9692 (
            .O(N__39280),
            .I(N__39224));
    LocalMux I__9691 (
            .O(N__39277),
            .I(N__39224));
    Span4Mux_h I__9690 (
            .O(N__39272),
            .I(N__39221));
    InMux I__9689 (
            .O(N__39271),
            .I(N__39216));
    InMux I__9688 (
            .O(N__39270),
            .I(N__39216));
    InMux I__9687 (
            .O(N__39269),
            .I(N__39213));
    LocalMux I__9686 (
            .O(N__39266),
            .I(N__39210));
    LocalMux I__9685 (
            .O(N__39263),
            .I(N__39193));
    LocalMux I__9684 (
            .O(N__39258),
            .I(N__39193));
    LocalMux I__9683 (
            .O(N__39255),
            .I(N__39193));
    LocalMux I__9682 (
            .O(N__39252),
            .I(N__39193));
    LocalMux I__9681 (
            .O(N__39247),
            .I(N__39193));
    Sp12to4 I__9680 (
            .O(N__39244),
            .I(N__39193));
    LocalMux I__9679 (
            .O(N__39241),
            .I(N__39193));
    LocalMux I__9678 (
            .O(N__39238),
            .I(N__39193));
    Span4Mux_v I__9677 (
            .O(N__39231),
            .I(N__39190));
    Span4Mux_v I__9676 (
            .O(N__39224),
            .I(N__39187));
    Sp12to4 I__9675 (
            .O(N__39221),
            .I(N__39178));
    LocalMux I__9674 (
            .O(N__39216),
            .I(N__39178));
    LocalMux I__9673 (
            .O(N__39213),
            .I(N__39178));
    Span12Mux_h I__9672 (
            .O(N__39210),
            .I(N__39178));
    Span12Mux_v I__9671 (
            .O(N__39193),
            .I(N__39175));
    Span4Mux_h I__9670 (
            .O(N__39190),
            .I(N__39172));
    Odrv4 I__9669 (
            .O(N__39187),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv12 I__9668 (
            .O(N__39178),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv12 I__9667 (
            .O(N__39175),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__9666 (
            .O(N__39172),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    InMux I__9665 (
            .O(N__39163),
            .I(N__39160));
    LocalMux I__9664 (
            .O(N__39160),
            .I(N__39157));
    Odrv4 I__9663 (
            .O(N__39157),
            .I(N_436));
    InMux I__9662 (
            .O(N__39154),
            .I(N__39151));
    LocalMux I__9661 (
            .O(N__39151),
            .I(M_this_oam_ram_read_data_30));
    InMux I__9660 (
            .O(N__39148),
            .I(N__39145));
    LocalMux I__9659 (
            .O(N__39145),
            .I(N__39142));
    Span4Mux_h I__9658 (
            .O(N__39142),
            .I(N__39139));
    Span4Mux_h I__9657 (
            .O(N__39139),
            .I(N__39136));
    Odrv4 I__9656 (
            .O(N__39136),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_30 ));
    InMux I__9655 (
            .O(N__39133),
            .I(N__39130));
    LocalMux I__9654 (
            .O(N__39130),
            .I(N__39127));
    Span4Mux_h I__9653 (
            .O(N__39127),
            .I(N__39124));
    Odrv4 I__9652 (
            .O(N__39124),
            .I(M_this_oam_ram_read_data_9));
    InMux I__9651 (
            .O(N__39121),
            .I(N__39118));
    LocalMux I__9650 (
            .O(N__39118),
            .I(N__39115));
    Span4Mux_v I__9649 (
            .O(N__39115),
            .I(N__39112));
    Odrv4 I__9648 (
            .O(N__39112),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_9 ));
    InMux I__9647 (
            .O(N__39109),
            .I(N__39106));
    LocalMux I__9646 (
            .O(N__39106),
            .I(N_435));
    InMux I__9645 (
            .O(N__39103),
            .I(N__39099));
    InMux I__9644 (
            .O(N__39102),
            .I(N__39096));
    LocalMux I__9643 (
            .O(N__39099),
            .I(N__39093));
    LocalMux I__9642 (
            .O(N__39096),
            .I(N__39087));
    Span4Mux_h I__9641 (
            .O(N__39093),
            .I(N__39087));
    InMux I__9640 (
            .O(N__39092),
            .I(N__39084));
    Span4Mux_v I__9639 (
            .O(N__39087),
            .I(N__39078));
    LocalMux I__9638 (
            .O(N__39084),
            .I(N__39075));
    InMux I__9637 (
            .O(N__39083),
            .I(N__39068));
    InMux I__9636 (
            .O(N__39082),
            .I(N__39068));
    InMux I__9635 (
            .O(N__39081),
            .I(N__39068));
    Odrv4 I__9634 (
            .O(N__39078),
            .I(M_this_oam_ram_read_data_17));
    Odrv4 I__9633 (
            .O(N__39075),
            .I(M_this_oam_ram_read_data_17));
    LocalMux I__9632 (
            .O(N__39068),
            .I(M_this_oam_ram_read_data_17));
    InMux I__9631 (
            .O(N__39061),
            .I(N__39058));
    LocalMux I__9630 (
            .O(N__39058),
            .I(N__39053));
    InMux I__9629 (
            .O(N__39057),
            .I(N__39050));
    InMux I__9628 (
            .O(N__39056),
            .I(N__39047));
    Sp12to4 I__9627 (
            .O(N__39053),
            .I(N__39041));
    LocalMux I__9626 (
            .O(N__39050),
            .I(N__39041));
    LocalMux I__9625 (
            .O(N__39047),
            .I(N__39038));
    InMux I__9624 (
            .O(N__39046),
            .I(N__39035));
    Span12Mux_v I__9623 (
            .O(N__39041),
            .I(N__39029));
    Span4Mux_v I__9622 (
            .O(N__39038),
            .I(N__39024));
    LocalMux I__9621 (
            .O(N__39035),
            .I(N__39024));
    InMux I__9620 (
            .O(N__39034),
            .I(N__39017));
    InMux I__9619 (
            .O(N__39033),
            .I(N__39017));
    InMux I__9618 (
            .O(N__39032),
            .I(N__39017));
    Odrv12 I__9617 (
            .O(N__39029),
            .I(M_this_oam_ram_read_data_16));
    Odrv4 I__9616 (
            .O(N__39024),
            .I(M_this_oam_ram_read_data_16));
    LocalMux I__9615 (
            .O(N__39017),
            .I(M_this_oam_ram_read_data_16));
    InMux I__9614 (
            .O(N__39010),
            .I(N__39007));
    LocalMux I__9613 (
            .O(N__39007),
            .I(N__39004));
    Span12Mux_v I__9612 (
            .O(N__39004),
            .I(N__39001));
    Odrv12 I__9611 (
            .O(N__39001),
            .I(\this_ppu.un1_oam_data_1_1 ));
    InMux I__9610 (
            .O(N__38998),
            .I(N__38995));
    LocalMux I__9609 (
            .O(N__38995),
            .I(\this_spr_ram.mem_out_bus5_2 ));
    InMux I__9608 (
            .O(N__38992),
            .I(N__38989));
    LocalMux I__9607 (
            .O(N__38989),
            .I(N__38986));
    Span4Mux_v I__9606 (
            .O(N__38986),
            .I(N__38983));
    Odrv4 I__9605 (
            .O(N__38983),
            .I(\this_spr_ram.mem_out_bus1_2 ));
    InMux I__9604 (
            .O(N__38980),
            .I(N__38977));
    LocalMux I__9603 (
            .O(N__38977),
            .I(N__38974));
    Span4Mux_h I__9602 (
            .O(N__38974),
            .I(N__38971));
    Sp12to4 I__9601 (
            .O(N__38971),
            .I(N__38968));
    Odrv12 I__9600 (
            .O(N__38968),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ));
    InMux I__9599 (
            .O(N__38965),
            .I(N__38962));
    LocalMux I__9598 (
            .O(N__38962),
            .I(N__38959));
    Odrv4 I__9597 (
            .O(N__38959),
            .I(\this_spr_ram.mem_out_bus5_0 ));
    InMux I__9596 (
            .O(N__38956),
            .I(N__38953));
    LocalMux I__9595 (
            .O(N__38953),
            .I(N__38950));
    Span4Mux_v I__9594 (
            .O(N__38950),
            .I(N__38947));
    Odrv4 I__9593 (
            .O(N__38947),
            .I(\this_spr_ram.mem_out_bus1_0 ));
    InMux I__9592 (
            .O(N__38944),
            .I(N__38938));
    InMux I__9591 (
            .O(N__38943),
            .I(N__38938));
    LocalMux I__9590 (
            .O(N__38938),
            .I(N__38925));
    InMux I__9589 (
            .O(N__38937),
            .I(N__38920));
    InMux I__9588 (
            .O(N__38936),
            .I(N__38920));
    InMux I__9587 (
            .O(N__38935),
            .I(N__38915));
    InMux I__9586 (
            .O(N__38934),
            .I(N__38915));
    InMux I__9585 (
            .O(N__38933),
            .I(N__38911));
    InMux I__9584 (
            .O(N__38932),
            .I(N__38908));
    InMux I__9583 (
            .O(N__38931),
            .I(N__38905));
    InMux I__9582 (
            .O(N__38930),
            .I(N__38902));
    InMux I__9581 (
            .O(N__38929),
            .I(N__38896));
    InMux I__9580 (
            .O(N__38928),
            .I(N__38893));
    Span4Mux_v I__9579 (
            .O(N__38925),
            .I(N__38886));
    LocalMux I__9578 (
            .O(N__38920),
            .I(N__38886));
    LocalMux I__9577 (
            .O(N__38915),
            .I(N__38886));
    InMux I__9576 (
            .O(N__38914),
            .I(N__38883));
    LocalMux I__9575 (
            .O(N__38911),
            .I(N__38880));
    LocalMux I__9574 (
            .O(N__38908),
            .I(N__38873));
    LocalMux I__9573 (
            .O(N__38905),
            .I(N__38873));
    LocalMux I__9572 (
            .O(N__38902),
            .I(N__38873));
    InMux I__9571 (
            .O(N__38901),
            .I(N__38870));
    InMux I__9570 (
            .O(N__38900),
            .I(N__38867));
    InMux I__9569 (
            .O(N__38899),
            .I(N__38864));
    LocalMux I__9568 (
            .O(N__38896),
            .I(N__38859));
    LocalMux I__9567 (
            .O(N__38893),
            .I(N__38859));
    Span4Mux_h I__9566 (
            .O(N__38886),
            .I(N__38856));
    LocalMux I__9565 (
            .O(N__38883),
            .I(N__38853));
    Span4Mux_h I__9564 (
            .O(N__38880),
            .I(N__38848));
    Span4Mux_v I__9563 (
            .O(N__38873),
            .I(N__38848));
    LocalMux I__9562 (
            .O(N__38870),
            .I(N__38845));
    LocalMux I__9561 (
            .O(N__38867),
            .I(N__38842));
    LocalMux I__9560 (
            .O(N__38864),
            .I(N__38837));
    Span4Mux_v I__9559 (
            .O(N__38859),
            .I(N__38837));
    Span4Mux_h I__9558 (
            .O(N__38856),
            .I(N__38834));
    Span12Mux_h I__9557 (
            .O(N__38853),
            .I(N__38831));
    Span4Mux_h I__9556 (
            .O(N__38848),
            .I(N__38828));
    Span12Mux_h I__9555 (
            .O(N__38845),
            .I(N__38825));
    Odrv4 I__9554 (
            .O(N__38842),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__9553 (
            .O(N__38837),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__9552 (
            .O(N__38834),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv12 I__9551 (
            .O(N__38831),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__9550 (
            .O(N__38828),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv12 I__9549 (
            .O(N__38825),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    InMux I__9548 (
            .O(N__38812),
            .I(N__38809));
    LocalMux I__9547 (
            .O(N__38809),
            .I(N__38806));
    Span12Mux_h I__9546 (
            .O(N__38806),
            .I(N__38803));
    Odrv12 I__9545 (
            .O(N__38803),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ));
    InMux I__9544 (
            .O(N__38800),
            .I(N__38797));
    LocalMux I__9543 (
            .O(N__38797),
            .I(N__38794));
    Odrv4 I__9542 (
            .O(N__38794),
            .I(un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0));
    InMux I__9541 (
            .O(N__38791),
            .I(N__38788));
    LocalMux I__9540 (
            .O(N__38788),
            .I(N__38785));
    Span4Mux_v I__9539 (
            .O(N__38785),
            .I(N__38781));
    InMux I__9538 (
            .O(N__38784),
            .I(N__38776));
    Span4Mux_v I__9537 (
            .O(N__38781),
            .I(N__38773));
    InMux I__9536 (
            .O(N__38780),
            .I(N__38770));
    InMux I__9535 (
            .O(N__38779),
            .I(N__38766));
    LocalMux I__9534 (
            .O(N__38776),
            .I(N__38761));
    Span4Mux_v I__9533 (
            .O(N__38773),
            .I(N__38755));
    LocalMux I__9532 (
            .O(N__38770),
            .I(N__38755));
    InMux I__9531 (
            .O(N__38769),
            .I(N__38751));
    LocalMux I__9530 (
            .O(N__38766),
            .I(N__38748));
    InMux I__9529 (
            .O(N__38765),
            .I(N__38745));
    InMux I__9528 (
            .O(N__38764),
            .I(N__38742));
    Span4Mux_v I__9527 (
            .O(N__38761),
            .I(N__38739));
    CascadeMux I__9526 (
            .O(N__38760),
            .I(N__38736));
    Span4Mux_v I__9525 (
            .O(N__38755),
            .I(N__38733));
    InMux I__9524 (
            .O(N__38754),
            .I(N__38730));
    LocalMux I__9523 (
            .O(N__38751),
            .I(N__38727));
    Span4Mux_h I__9522 (
            .O(N__38748),
            .I(N__38722));
    LocalMux I__9521 (
            .O(N__38745),
            .I(N__38722));
    LocalMux I__9520 (
            .O(N__38742),
            .I(N__38719));
    Span4Mux_h I__9519 (
            .O(N__38739),
            .I(N__38716));
    InMux I__9518 (
            .O(N__38736),
            .I(N__38713));
    Span4Mux_h I__9517 (
            .O(N__38733),
            .I(N__38710));
    LocalMux I__9516 (
            .O(N__38730),
            .I(N__38707));
    Span12Mux_v I__9515 (
            .O(N__38727),
            .I(N__38704));
    Span4Mux_v I__9514 (
            .O(N__38722),
            .I(N__38701));
    Span12Mux_h I__9513 (
            .O(N__38719),
            .I(N__38698));
    Span4Mux_h I__9512 (
            .O(N__38716),
            .I(N__38693));
    LocalMux I__9511 (
            .O(N__38713),
            .I(N__38693));
    Span4Mux_h I__9510 (
            .O(N__38710),
            .I(N__38688));
    Span4Mux_v I__9509 (
            .O(N__38707),
            .I(N__38688));
    Span12Mux_h I__9508 (
            .O(N__38704),
            .I(N__38685));
    Span4Mux_h I__9507 (
            .O(N__38701),
            .I(N__38682));
    Span12Mux_h I__9506 (
            .O(N__38698),
            .I(N__38677));
    Sp12to4 I__9505 (
            .O(N__38693),
            .I(N__38677));
    IoSpan4Mux I__9504 (
            .O(N__38688),
            .I(N__38674));
    Odrv12 I__9503 (
            .O(N__38685),
            .I(port_data_c_2));
    Odrv4 I__9502 (
            .O(N__38682),
            .I(port_data_c_2));
    Odrv12 I__9501 (
            .O(N__38677),
            .I(port_data_c_2));
    Odrv4 I__9500 (
            .O(N__38674),
            .I(port_data_c_2));
    IoInMux I__9499 (
            .O(N__38665),
            .I(N__38662));
    LocalMux I__9498 (
            .O(N__38662),
            .I(N__38659));
    IoSpan4Mux I__9497 (
            .O(N__38659),
            .I(N__38656));
    Span4Mux_s2_v I__9496 (
            .O(N__38656),
            .I(N__38653));
    Sp12to4 I__9495 (
            .O(N__38653),
            .I(N__38649));
    InMux I__9494 (
            .O(N__38652),
            .I(N__38646));
    Span12Mux_s10_v I__9493 (
            .O(N__38649),
            .I(N__38641));
    LocalMux I__9492 (
            .O(N__38646),
            .I(N__38641));
    Odrv12 I__9491 (
            .O(N__38641),
            .I(M_this_ext_address_qZ0Z_10));
    InMux I__9490 (
            .O(N__38638),
            .I(N__38635));
    LocalMux I__9489 (
            .O(N__38635),
            .I(N__38632));
    Span4Mux_v I__9488 (
            .O(N__38632),
            .I(N__38629));
    Odrv4 I__9487 (
            .O(N__38629),
            .I(un1_M_this_ext_address_q_cry_3_THRU_CO));
    IoInMux I__9486 (
            .O(N__38626),
            .I(N__38622));
    InMux I__9485 (
            .O(N__38625),
            .I(N__38619));
    LocalMux I__9484 (
            .O(N__38622),
            .I(N__38616));
    LocalMux I__9483 (
            .O(N__38619),
            .I(N__38612));
    Span12Mux_s6_h I__9482 (
            .O(N__38616),
            .I(N__38609));
    InMux I__9481 (
            .O(N__38615),
            .I(N__38606));
    Span4Mux_v I__9480 (
            .O(N__38612),
            .I(N__38603));
    Odrv12 I__9479 (
            .O(N__38609),
            .I(M_this_ext_address_qZ0Z_4));
    LocalMux I__9478 (
            .O(N__38606),
            .I(M_this_ext_address_qZ0Z_4));
    Odrv4 I__9477 (
            .O(N__38603),
            .I(M_this_ext_address_qZ0Z_4));
    InMux I__9476 (
            .O(N__38596),
            .I(N__38593));
    LocalMux I__9475 (
            .O(N__38593),
            .I(N__38590));
    Span4Mux_v I__9474 (
            .O(N__38590),
            .I(N__38587));
    Span4Mux_h I__9473 (
            .O(N__38587),
            .I(N__38584));
    Odrv4 I__9472 (
            .O(N__38584),
            .I(\this_ppu.un1_oam_data_1_4 ));
    InMux I__9471 (
            .O(N__38581),
            .I(N__38578));
    LocalMux I__9470 (
            .O(N__38578),
            .I(M_this_oam_ram_read_data_31));
    InMux I__9469 (
            .O(N__38575),
            .I(N__38572));
    LocalMux I__9468 (
            .O(N__38572),
            .I(N__38569));
    Odrv4 I__9467 (
            .O(N__38569),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_31 ));
    InMux I__9466 (
            .O(N__38566),
            .I(N__38560));
    InMux I__9465 (
            .O(N__38565),
            .I(N__38557));
    CascadeMux I__9464 (
            .O(N__38564),
            .I(N__38553));
    CascadeMux I__9463 (
            .O(N__38563),
            .I(N__38550));
    LocalMux I__9462 (
            .O(N__38560),
            .I(N__38547));
    LocalMux I__9461 (
            .O(N__38557),
            .I(N__38544));
    InMux I__9460 (
            .O(N__38556),
            .I(N__38537));
    InMux I__9459 (
            .O(N__38553),
            .I(N__38537));
    InMux I__9458 (
            .O(N__38550),
            .I(N__38537));
    Span4Mux_v I__9457 (
            .O(N__38547),
            .I(N__38534));
    Span4Mux_h I__9456 (
            .O(N__38544),
            .I(N__38529));
    LocalMux I__9455 (
            .O(N__38537),
            .I(N__38529));
    Span4Mux_v I__9454 (
            .O(N__38534),
            .I(N__38526));
    Odrv4 I__9453 (
            .O(N__38529),
            .I(M_this_oam_ram_read_data_19));
    Odrv4 I__9452 (
            .O(N__38526),
            .I(M_this_oam_ram_read_data_19));
    InMux I__9451 (
            .O(N__38521),
            .I(N__38518));
    LocalMux I__9450 (
            .O(N__38518),
            .I(N__38515));
    Odrv4 I__9449 (
            .O(N__38515),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_19 ));
    CascadeMux I__9448 (
            .O(N__38512),
            .I(N__38509));
    InMux I__9447 (
            .O(N__38509),
            .I(N__38505));
    InMux I__9446 (
            .O(N__38508),
            .I(N__38502));
    LocalMux I__9445 (
            .O(N__38505),
            .I(N__38497));
    LocalMux I__9444 (
            .O(N__38502),
            .I(N__38494));
    InMux I__9443 (
            .O(N__38501),
            .I(N__38489));
    InMux I__9442 (
            .O(N__38500),
            .I(N__38489));
    Span4Mux_h I__9441 (
            .O(N__38497),
            .I(N__38486));
    Span4Mux_h I__9440 (
            .O(N__38494),
            .I(N__38481));
    LocalMux I__9439 (
            .O(N__38489),
            .I(N__38481));
    Span4Mux_v I__9438 (
            .O(N__38486),
            .I(N__38478));
    Odrv4 I__9437 (
            .O(N__38481),
            .I(M_this_oam_ram_read_data_20));
    Odrv4 I__9436 (
            .O(N__38478),
            .I(M_this_oam_ram_read_data_20));
    InMux I__9435 (
            .O(N__38473),
            .I(N__38470));
    LocalMux I__9434 (
            .O(N__38470),
            .I(N__38467));
    Span4Mux_h I__9433 (
            .O(N__38467),
            .I(N__38464));
    Odrv4 I__9432 (
            .O(N__38464),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_20 ));
    InMux I__9431 (
            .O(N__38461),
            .I(N__38458));
    LocalMux I__9430 (
            .O(N__38458),
            .I(M_this_oam_ram_read_data_24));
    InMux I__9429 (
            .O(N__38455),
            .I(N__38452));
    LocalMux I__9428 (
            .O(N__38452),
            .I(N__38449));
    Span4Mux_h I__9427 (
            .O(N__38449),
            .I(N__38446));
    Odrv4 I__9426 (
            .O(N__38446),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_24 ));
    InMux I__9425 (
            .O(N__38443),
            .I(N__38438));
    InMux I__9424 (
            .O(N__38442),
            .I(N__38435));
    InMux I__9423 (
            .O(N__38441),
            .I(N__38432));
    LocalMux I__9422 (
            .O(N__38438),
            .I(N__38427));
    LocalMux I__9421 (
            .O(N__38435),
            .I(N__38424));
    LocalMux I__9420 (
            .O(N__38432),
            .I(N__38421));
    InMux I__9419 (
            .O(N__38431),
            .I(N__38416));
    InMux I__9418 (
            .O(N__38430),
            .I(N__38416));
    Span4Mux_v I__9417 (
            .O(N__38427),
            .I(N__38412));
    Span12Mux_v I__9416 (
            .O(N__38424),
            .I(N__38409));
    Span4Mux_h I__9415 (
            .O(N__38421),
            .I(N__38404));
    LocalMux I__9414 (
            .O(N__38416),
            .I(N__38404));
    InMux I__9413 (
            .O(N__38415),
            .I(N__38401));
    Span4Mux_v I__9412 (
            .O(N__38412),
            .I(N__38398));
    Odrv12 I__9411 (
            .O(N__38409),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__9410 (
            .O(N__38404),
            .I(M_this_oam_ram_read_data_18));
    LocalMux I__9409 (
            .O(N__38401),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__9408 (
            .O(N__38398),
            .I(M_this_oam_ram_read_data_18));
    InMux I__9407 (
            .O(N__38389),
            .I(N__38386));
    LocalMux I__9406 (
            .O(N__38386),
            .I(N__38383));
    Span4Mux_h I__9405 (
            .O(N__38383),
            .I(N__38380));
    Span4Mux_v I__9404 (
            .O(N__38380),
            .I(N__38377));
    Odrv4 I__9403 (
            .O(N__38377),
            .I(\this_ppu.un1_oam_data_1_2 ));
    InMux I__9402 (
            .O(N__38374),
            .I(N__38371));
    LocalMux I__9401 (
            .O(N__38371),
            .I(N__38368));
    Odrv12 I__9400 (
            .O(N__38368),
            .I(M_this_data_tmp_qZ0Z_17));
    InMux I__9399 (
            .O(N__38365),
            .I(N__38362));
    LocalMux I__9398 (
            .O(N__38362),
            .I(M_this_oam_ram_write_data_17));
    InMux I__9397 (
            .O(N__38359),
            .I(N__38356));
    LocalMux I__9396 (
            .O(N__38356),
            .I(N__38352));
    InMux I__9395 (
            .O(N__38355),
            .I(N__38349));
    Span4Mux_v I__9394 (
            .O(N__38352),
            .I(N__38346));
    LocalMux I__9393 (
            .O(N__38349),
            .I(\this_ppu.un1_oam_data_1_4_c2 ));
    Odrv4 I__9392 (
            .O(N__38346),
            .I(\this_ppu.un1_oam_data_1_4_c2 ));
    InMux I__9391 (
            .O(N__38341),
            .I(N__38335));
    InMux I__9390 (
            .O(N__38340),
            .I(N__38335));
    LocalMux I__9389 (
            .O(N__38335),
            .I(M_this_oam_ram_read_data_5));
    InMux I__9388 (
            .O(N__38332),
            .I(N__38329));
    LocalMux I__9387 (
            .O(N__38329),
            .I(N__38326));
    Span4Mux_h I__9386 (
            .O(N__38326),
            .I(N__38323));
    Odrv4 I__9385 (
            .O(N__38323),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_5 ));
    InMux I__9384 (
            .O(N__38320),
            .I(N__38314));
    InMux I__9383 (
            .O(N__38319),
            .I(N__38314));
    LocalMux I__9382 (
            .O(N__38314),
            .I(M_this_oam_ram_read_data_6));
    InMux I__9381 (
            .O(N__38311),
            .I(N__38308));
    LocalMux I__9380 (
            .O(N__38308),
            .I(N__38305));
    Odrv4 I__9379 (
            .O(N__38305),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_6 ));
    CascadeMux I__9378 (
            .O(N__38302),
            .I(N__38298));
    InMux I__9377 (
            .O(N__38301),
            .I(N__38293));
    InMux I__9376 (
            .O(N__38298),
            .I(N__38293));
    LocalMux I__9375 (
            .O(N__38293),
            .I(M_this_oam_ram_read_data_7));
    InMux I__9374 (
            .O(N__38290),
            .I(N__38287));
    LocalMux I__9373 (
            .O(N__38287),
            .I(N__38284));
    Odrv4 I__9372 (
            .O(N__38284),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_7 ));
    InMux I__9371 (
            .O(N__38281),
            .I(N__38278));
    LocalMux I__9370 (
            .O(N__38278),
            .I(N__38275));
    Odrv4 I__9369 (
            .O(N__38275),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_0 ));
    InMux I__9368 (
            .O(N__38272),
            .I(N__38269));
    LocalMux I__9367 (
            .O(N__38269),
            .I(N__38266));
    Span4Mux_h I__9366 (
            .O(N__38266),
            .I(N__38263));
    Odrv4 I__9365 (
            .O(N__38263),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_1 ));
    InMux I__9364 (
            .O(N__38260),
            .I(N__38257));
    LocalMux I__9363 (
            .O(N__38257),
            .I(N__38253));
    InMux I__9362 (
            .O(N__38256),
            .I(N__38250));
    Odrv4 I__9361 (
            .O(N__38253),
            .I(M_this_oam_ram_read_data_2));
    LocalMux I__9360 (
            .O(N__38250),
            .I(M_this_oam_ram_read_data_2));
    InMux I__9359 (
            .O(N__38245),
            .I(N__38239));
    InMux I__9358 (
            .O(N__38244),
            .I(N__38239));
    LocalMux I__9357 (
            .O(N__38239),
            .I(M_this_oam_ram_read_data_1));
    InMux I__9356 (
            .O(N__38236),
            .I(N__38232));
    CascadeMux I__9355 (
            .O(N__38235),
            .I(N__38229));
    LocalMux I__9354 (
            .O(N__38232),
            .I(N__38226));
    InMux I__9353 (
            .O(N__38229),
            .I(N__38223));
    Odrv4 I__9352 (
            .O(N__38226),
            .I(M_this_oam_ram_read_data_3));
    LocalMux I__9351 (
            .O(N__38223),
            .I(M_this_oam_ram_read_data_3));
    InMux I__9350 (
            .O(N__38218),
            .I(N__38212));
    InMux I__9349 (
            .O(N__38217),
            .I(N__38212));
    LocalMux I__9348 (
            .O(N__38212),
            .I(M_this_oam_ram_read_data_0));
    InMux I__9347 (
            .O(N__38209),
            .I(N__38206));
    LocalMux I__9346 (
            .O(N__38206),
            .I(N__38203));
    Odrv4 I__9345 (
            .O(N__38203),
            .I(\this_ppu.un12lto7Z0Z_5 ));
    InMux I__9344 (
            .O(N__38200),
            .I(N__38197));
    LocalMux I__9343 (
            .O(N__38197),
            .I(M_this_oam_ram_read_data_27));
    InMux I__9342 (
            .O(N__38194),
            .I(N__38191));
    LocalMux I__9341 (
            .O(N__38191),
            .I(N__38188));
    Span4Mux_h I__9340 (
            .O(N__38188),
            .I(N__38185));
    Odrv4 I__9339 (
            .O(N__38185),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_27 ));
    InMux I__9338 (
            .O(N__38182),
            .I(N__38179));
    LocalMux I__9337 (
            .O(N__38179),
            .I(N__38176));
    Span4Mux_h I__9336 (
            .O(N__38176),
            .I(N__38173));
    Span4Mux_v I__9335 (
            .O(N__38173),
            .I(N__38170));
    Odrv4 I__9334 (
            .O(N__38170),
            .I(\this_ppu.un1_oam_data_1_3 ));
    InMux I__9333 (
            .O(N__38167),
            .I(N__38164));
    LocalMux I__9332 (
            .O(N__38164),
            .I(M_this_oam_ram_read_data_29));
    InMux I__9331 (
            .O(N__38161),
            .I(N__38158));
    LocalMux I__9330 (
            .O(N__38158),
            .I(N__38155));
    Span4Mux_h I__9329 (
            .O(N__38155),
            .I(N__38152));
    Odrv4 I__9328 (
            .O(N__38152),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_29 ));
    InMux I__9327 (
            .O(N__38149),
            .I(N__38146));
    LocalMux I__9326 (
            .O(N__38146),
            .I(N__38143));
    Span4Mux_h I__9325 (
            .O(N__38143),
            .I(N__38140));
    Odrv4 I__9324 (
            .O(N__38140),
            .I(M_this_oam_ram_read_data_25));
    InMux I__9323 (
            .O(N__38137),
            .I(N__38134));
    LocalMux I__9322 (
            .O(N__38134),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_25 ));
    InMux I__9321 (
            .O(N__38131),
            .I(N__38128));
    LocalMux I__9320 (
            .O(N__38128),
            .I(N__38125));
    Span4Mux_v I__9319 (
            .O(N__38125),
            .I(N__38122));
    Odrv4 I__9318 (
            .O(N__38122),
            .I(M_this_oam_ram_read_data_26));
    InMux I__9317 (
            .O(N__38119),
            .I(N__38116));
    LocalMux I__9316 (
            .O(N__38116),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_26 ));
    InMux I__9315 (
            .O(N__38113),
            .I(N__38110));
    LocalMux I__9314 (
            .O(N__38110),
            .I(N__38107));
    Span12Mux_s9_h I__9313 (
            .O(N__38107),
            .I(N__38104));
    Odrv12 I__9312 (
            .O(N__38104),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__9311 (
            .O(N__38101),
            .I(N__38098));
    LocalMux I__9310 (
            .O(N__38098),
            .I(M_this_oam_ram_write_data_10));
    InMux I__9309 (
            .O(N__38095),
            .I(N__38092));
    LocalMux I__9308 (
            .O(N__38092),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__9307 (
            .O(N__38089),
            .I(N__38086));
    LocalMux I__9306 (
            .O(N__38086),
            .I(N__38083));
    Odrv4 I__9305 (
            .O(N__38083),
            .I(M_this_oam_ram_write_data_6));
    InMux I__9304 (
            .O(N__38080),
            .I(N__38077));
    LocalMux I__9303 (
            .O(N__38077),
            .I(N__38074));
    Span4Mux_h I__9302 (
            .O(N__38074),
            .I(N__38071));
    Span4Mux_h I__9301 (
            .O(N__38071),
            .I(N__38068));
    Odrv4 I__9300 (
            .O(N__38068),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__9299 (
            .O(N__38065),
            .I(N__38062));
    LocalMux I__9298 (
            .O(N__38062),
            .I(N__38059));
    Odrv4 I__9297 (
            .O(N__38059),
            .I(M_this_oam_ram_write_data_11));
    InMux I__9296 (
            .O(N__38056),
            .I(N__38053));
    LocalMux I__9295 (
            .O(N__38053),
            .I(N__38050));
    Span4Mux_h I__9294 (
            .O(N__38050),
            .I(N__38047));
    Odrv4 I__9293 (
            .O(N__38047),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_2 ));
    InMux I__9292 (
            .O(N__38044),
            .I(N__38041));
    LocalMux I__9291 (
            .O(N__38041),
            .I(N__38038));
    Odrv4 I__9290 (
            .O(N__38038),
            .I(\this_ppu.un12lto7Z0Z_4 ));
    InMux I__9289 (
            .O(N__38035),
            .I(N__38029));
    InMux I__9288 (
            .O(N__38034),
            .I(N__38029));
    LocalMux I__9287 (
            .O(N__38029),
            .I(M_this_oam_ram_read_data_4));
    InMux I__9286 (
            .O(N__38026),
            .I(N__38023));
    LocalMux I__9285 (
            .O(N__38023),
            .I(N__38020));
    Span4Mux_h I__9284 (
            .O(N__38020),
            .I(N__38017));
    Odrv4 I__9283 (
            .O(N__38017),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_4 ));
    InMux I__9282 (
            .O(N__38014),
            .I(un1_M_this_ext_address_q_cry_12));
    IoInMux I__9281 (
            .O(N__38011),
            .I(N__38008));
    LocalMux I__9280 (
            .O(N__38008),
            .I(N__38005));
    Span4Mux_s1_h I__9279 (
            .O(N__38005),
            .I(N__38002));
    Sp12to4 I__9278 (
            .O(N__38002),
            .I(N__37998));
    CascadeMux I__9277 (
            .O(N__38001),
            .I(N__37995));
    Span12Mux_v I__9276 (
            .O(N__37998),
            .I(N__37992));
    InMux I__9275 (
            .O(N__37995),
            .I(N__37989));
    Odrv12 I__9274 (
            .O(N__37992),
            .I(M_this_ext_address_qZ0Z_14));
    LocalMux I__9273 (
            .O(N__37989),
            .I(M_this_ext_address_qZ0Z_14));
    InMux I__9272 (
            .O(N__37984),
            .I(N__37981));
    LocalMux I__9271 (
            .O(N__37981),
            .I(un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0));
    InMux I__9270 (
            .O(N__37978),
            .I(un1_M_this_ext_address_q_cry_13));
    IoInMux I__9269 (
            .O(N__37975),
            .I(N__37972));
    LocalMux I__9268 (
            .O(N__37972),
            .I(N__37969));
    Span4Mux_s0_h I__9267 (
            .O(N__37969),
            .I(N__37966));
    Sp12to4 I__9266 (
            .O(N__37966),
            .I(N__37962));
    InMux I__9265 (
            .O(N__37965),
            .I(N__37959));
    Span12Mux_v I__9264 (
            .O(N__37962),
            .I(N__37956));
    LocalMux I__9263 (
            .O(N__37959),
            .I(N__37953));
    Odrv12 I__9262 (
            .O(N__37956),
            .I(M_this_ext_address_qZ0Z_15));
    Odrv4 I__9261 (
            .O(N__37953),
            .I(M_this_ext_address_qZ0Z_15));
    InMux I__9260 (
            .O(N__37948),
            .I(un1_M_this_ext_address_q_cry_14));
    InMux I__9259 (
            .O(N__37945),
            .I(N__37942));
    LocalMux I__9258 (
            .O(N__37942),
            .I(N__37939));
    Odrv4 I__9257 (
            .O(N__37939),
            .I(un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0));
    InMux I__9256 (
            .O(N__37936),
            .I(N__37933));
    LocalMux I__9255 (
            .O(N__37933),
            .I(N__37930));
    Odrv4 I__9254 (
            .O(N__37930),
            .I(M_this_oam_ram_read_data_13));
    InMux I__9253 (
            .O(N__37927),
            .I(N__37924));
    LocalMux I__9252 (
            .O(N__37924),
            .I(N__37921));
    Odrv4 I__9251 (
            .O(N__37921),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_13 ));
    InMux I__9250 (
            .O(N__37918),
            .I(N__37915));
    LocalMux I__9249 (
            .O(N__37915),
            .I(N__37912));
    Odrv4 I__9248 (
            .O(N__37912),
            .I(M_this_oam_ram_read_data_15));
    InMux I__9247 (
            .O(N__37909),
            .I(N__37906));
    LocalMux I__9246 (
            .O(N__37906),
            .I(N__37903));
    Odrv4 I__9245 (
            .O(N__37903),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_15 ));
    InMux I__9244 (
            .O(N__37900),
            .I(N__37897));
    LocalMux I__9243 (
            .O(N__37897),
            .I(N__37894));
    Odrv4 I__9242 (
            .O(N__37894),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_3 ));
    InMux I__9241 (
            .O(N__37891),
            .I(N__37888));
    LocalMux I__9240 (
            .O(N__37888),
            .I(N__37885));
    Odrv4 I__9239 (
            .O(N__37885),
            .I(M_this_oam_ram_read_data_8));
    InMux I__9238 (
            .O(N__37882),
            .I(N__37879));
    LocalMux I__9237 (
            .O(N__37879),
            .I(N__37876));
    Odrv4 I__9236 (
            .O(N__37876),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_8 ));
    InMux I__9235 (
            .O(N__37873),
            .I(N__37870));
    LocalMux I__9234 (
            .O(N__37870),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_16 ));
    InMux I__9233 (
            .O(N__37867),
            .I(N__37864));
    LocalMux I__9232 (
            .O(N__37864),
            .I(N__37861));
    Odrv4 I__9231 (
            .O(N__37861),
            .I(M_this_oam_ram_read_data_10));
    InMux I__9230 (
            .O(N__37858),
            .I(N__37855));
    LocalMux I__9229 (
            .O(N__37855),
            .I(N__37852));
    Odrv4 I__9228 (
            .O(N__37852),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_10 ));
    InMux I__9227 (
            .O(N__37849),
            .I(un1_M_this_ext_address_q_cry_3));
    InMux I__9226 (
            .O(N__37846),
            .I(un1_M_this_ext_address_q_cry_4));
    InMux I__9225 (
            .O(N__37843),
            .I(un1_M_this_ext_address_q_cry_5));
    InMux I__9224 (
            .O(N__37840),
            .I(un1_M_this_ext_address_q_cry_6));
    IoInMux I__9223 (
            .O(N__37837),
            .I(N__37834));
    LocalMux I__9222 (
            .O(N__37834),
            .I(N__37831));
    IoSpan4Mux I__9221 (
            .O(N__37831),
            .I(N__37828));
    IoSpan4Mux I__9220 (
            .O(N__37828),
            .I(N__37825));
    Span4Mux_s2_v I__9219 (
            .O(N__37825),
            .I(N__37822));
    Sp12to4 I__9218 (
            .O(N__37822),
            .I(N__37818));
    InMux I__9217 (
            .O(N__37821),
            .I(N__37815));
    Odrv12 I__9216 (
            .O(N__37818),
            .I(M_this_ext_address_qZ0Z_8));
    LocalMux I__9215 (
            .O(N__37815),
            .I(M_this_ext_address_qZ0Z_8));
    InMux I__9214 (
            .O(N__37810),
            .I(N__37807));
    LocalMux I__9213 (
            .O(N__37807),
            .I(un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0));
    InMux I__9212 (
            .O(N__37804),
            .I(bfn_24_22_0_));
    IoInMux I__9211 (
            .O(N__37801),
            .I(N__37798));
    LocalMux I__9210 (
            .O(N__37798),
            .I(N__37795));
    IoSpan4Mux I__9209 (
            .O(N__37795),
            .I(N__37792));
    Span4Mux_s3_v I__9208 (
            .O(N__37792),
            .I(N__37789));
    Span4Mux_v I__9207 (
            .O(N__37789),
            .I(N__37785));
    InMux I__9206 (
            .O(N__37788),
            .I(N__37782));
    Odrv4 I__9205 (
            .O(N__37785),
            .I(M_this_ext_address_qZ0Z_9));
    LocalMux I__9204 (
            .O(N__37782),
            .I(M_this_ext_address_qZ0Z_9));
    CascadeMux I__9203 (
            .O(N__37777),
            .I(N__37774));
    InMux I__9202 (
            .O(N__37774),
            .I(N__37771));
    LocalMux I__9201 (
            .O(N__37771),
            .I(N__37768));
    Odrv4 I__9200 (
            .O(N__37768),
            .I(un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0));
    InMux I__9199 (
            .O(N__37765),
            .I(un1_M_this_ext_address_q_cry_8));
    InMux I__9198 (
            .O(N__37762),
            .I(un1_M_this_ext_address_q_cry_9));
    InMux I__9197 (
            .O(N__37759),
            .I(un1_M_this_ext_address_q_cry_10));
    InMux I__9196 (
            .O(N__37756),
            .I(un1_M_this_ext_address_q_cry_11));
    InMux I__9195 (
            .O(N__37753),
            .I(N__37750));
    LocalMux I__9194 (
            .O(N__37750),
            .I(N__37747));
    Span12Mux_v I__9193 (
            .O(N__37747),
            .I(N__37744));
    Span12Mux_h I__9192 (
            .O(N__37744),
            .I(N__37740));
    InMux I__9191 (
            .O(N__37743),
            .I(N__37737));
    Odrv12 I__9190 (
            .O(N__37740),
            .I(M_this_ctrl_flags_qZ0Z_7));
    LocalMux I__9189 (
            .O(N__37737),
            .I(M_this_ctrl_flags_qZ0Z_7));
    InMux I__9188 (
            .O(N__37732),
            .I(N__37728));
    InMux I__9187 (
            .O(N__37731),
            .I(N__37725));
    LocalMux I__9186 (
            .O(N__37728),
            .I(N__37722));
    LocalMux I__9185 (
            .O(N__37725),
            .I(N_312_0));
    Odrv4 I__9184 (
            .O(N__37722),
            .I(N_312_0));
    IoInMux I__9183 (
            .O(N__37717),
            .I(N__37714));
    LocalMux I__9182 (
            .O(N__37714),
            .I(N__37711));
    Span4Mux_s0_v I__9181 (
            .O(N__37711),
            .I(N__37708));
    Sp12to4 I__9180 (
            .O(N__37708),
            .I(N__37705));
    Span12Mux_h I__9179 (
            .O(N__37705),
            .I(N__37701));
    CascadeMux I__9178 (
            .O(N__37704),
            .I(N__37697));
    Span12Mux_v I__9177 (
            .O(N__37701),
            .I(N__37694));
    InMux I__9176 (
            .O(N__37700),
            .I(N__37691));
    InMux I__9175 (
            .O(N__37697),
            .I(N__37688));
    Odrv12 I__9174 (
            .O(N__37694),
            .I(M_this_ext_address_qZ0Z_0));
    LocalMux I__9173 (
            .O(N__37691),
            .I(M_this_ext_address_qZ0Z_0));
    LocalMux I__9172 (
            .O(N__37688),
            .I(M_this_ext_address_qZ0Z_0));
    IoInMux I__9171 (
            .O(N__37681),
            .I(N__37678));
    LocalMux I__9170 (
            .O(N__37678),
            .I(N__37675));
    IoSpan4Mux I__9169 (
            .O(N__37675),
            .I(N__37672));
    Sp12to4 I__9168 (
            .O(N__37672),
            .I(N__37669));
    Span12Mux_v I__9167 (
            .O(N__37669),
            .I(N__37664));
    InMux I__9166 (
            .O(N__37668),
            .I(N__37661));
    InMux I__9165 (
            .O(N__37667),
            .I(N__37658));
    Odrv12 I__9164 (
            .O(N__37664),
            .I(M_this_ext_address_qZ0Z_1));
    LocalMux I__9163 (
            .O(N__37661),
            .I(M_this_ext_address_qZ0Z_1));
    LocalMux I__9162 (
            .O(N__37658),
            .I(M_this_ext_address_qZ0Z_1));
    CascadeMux I__9161 (
            .O(N__37651),
            .I(N__37648));
    InMux I__9160 (
            .O(N__37648),
            .I(N__37645));
    LocalMux I__9159 (
            .O(N__37645),
            .I(N__37642));
    Odrv4 I__9158 (
            .O(N__37642),
            .I(un1_M_this_ext_address_q_cry_0_THRU_CO));
    InMux I__9157 (
            .O(N__37639),
            .I(un1_M_this_ext_address_q_cry_0));
    IoInMux I__9156 (
            .O(N__37636),
            .I(N__37633));
    LocalMux I__9155 (
            .O(N__37633),
            .I(N__37630));
    Span12Mux_s0_v I__9154 (
            .O(N__37630),
            .I(N__37627));
    Span12Mux_v I__9153 (
            .O(N__37627),
            .I(N__37622));
    InMux I__9152 (
            .O(N__37626),
            .I(N__37619));
    InMux I__9151 (
            .O(N__37625),
            .I(N__37616));
    Odrv12 I__9150 (
            .O(N__37622),
            .I(M_this_ext_address_qZ0Z_2));
    LocalMux I__9149 (
            .O(N__37619),
            .I(M_this_ext_address_qZ0Z_2));
    LocalMux I__9148 (
            .O(N__37616),
            .I(M_this_ext_address_qZ0Z_2));
    InMux I__9147 (
            .O(N__37609),
            .I(N__37606));
    LocalMux I__9146 (
            .O(N__37606),
            .I(un1_M_this_ext_address_q_cry_1_THRU_CO));
    InMux I__9145 (
            .O(N__37603),
            .I(un1_M_this_ext_address_q_cry_1));
    IoInMux I__9144 (
            .O(N__37600),
            .I(N__37597));
    LocalMux I__9143 (
            .O(N__37597),
            .I(N__37594));
    Span4Mux_s1_h I__9142 (
            .O(N__37594),
            .I(N__37591));
    Span4Mux_h I__9141 (
            .O(N__37591),
            .I(N__37588));
    Span4Mux_v I__9140 (
            .O(N__37588),
            .I(N__37585));
    Span4Mux_v I__9139 (
            .O(N__37585),
            .I(N__37580));
    InMux I__9138 (
            .O(N__37584),
            .I(N__37577));
    InMux I__9137 (
            .O(N__37583),
            .I(N__37574));
    Odrv4 I__9136 (
            .O(N__37580),
            .I(M_this_ext_address_qZ0Z_3));
    LocalMux I__9135 (
            .O(N__37577),
            .I(M_this_ext_address_qZ0Z_3));
    LocalMux I__9134 (
            .O(N__37574),
            .I(M_this_ext_address_qZ0Z_3));
    CascadeMux I__9133 (
            .O(N__37567),
            .I(N__37564));
    InMux I__9132 (
            .O(N__37564),
            .I(N__37561));
    LocalMux I__9131 (
            .O(N__37561),
            .I(un1_M_this_ext_address_q_cry_2_THRU_CO));
    InMux I__9130 (
            .O(N__37558),
            .I(un1_M_this_ext_address_q_cry_2));
    InMux I__9129 (
            .O(N__37555),
            .I(N__37552));
    LocalMux I__9128 (
            .O(N__37552),
            .I(N__37544));
    InMux I__9127 (
            .O(N__37551),
            .I(N__37541));
    InMux I__9126 (
            .O(N__37550),
            .I(N__37538));
    InMux I__9125 (
            .O(N__37549),
            .I(N__37535));
    InMux I__9124 (
            .O(N__37548),
            .I(N__37530));
    InMux I__9123 (
            .O(N__37547),
            .I(N__37530));
    Span4Mux_v I__9122 (
            .O(N__37544),
            .I(N__37522));
    LocalMux I__9121 (
            .O(N__37541),
            .I(N__37522));
    LocalMux I__9120 (
            .O(N__37538),
            .I(N__37522));
    LocalMux I__9119 (
            .O(N__37535),
            .I(N__37519));
    LocalMux I__9118 (
            .O(N__37530),
            .I(N__37516));
    InMux I__9117 (
            .O(N__37529),
            .I(N__37513));
    Span4Mux_h I__9116 (
            .O(N__37522),
            .I(N__37510));
    Span4Mux_h I__9115 (
            .O(N__37519),
            .I(N__37507));
    Span4Mux_h I__9114 (
            .O(N__37516),
            .I(N__37504));
    LocalMux I__9113 (
            .O(N__37513),
            .I(N__37501));
    Span4Mux_v I__9112 (
            .O(N__37510),
            .I(N__37497));
    Span4Mux_v I__9111 (
            .O(N__37507),
            .I(N__37492));
    Span4Mux_h I__9110 (
            .O(N__37504),
            .I(N__37492));
    Span4Mux_h I__9109 (
            .O(N__37501),
            .I(N__37489));
    InMux I__9108 (
            .O(N__37500),
            .I(N__37486));
    Odrv4 I__9107 (
            .O(N__37497),
            .I(N_260_0));
    Odrv4 I__9106 (
            .O(N__37492),
            .I(N_260_0));
    Odrv4 I__9105 (
            .O(N__37489),
            .I(N_260_0));
    LocalMux I__9104 (
            .O(N__37486),
            .I(N_260_0));
    CascadeMux I__9103 (
            .O(N__37477),
            .I(N__37471));
    InMux I__9102 (
            .O(N__37476),
            .I(N__37468));
    CascadeMux I__9101 (
            .O(N__37475),
            .I(N__37463));
    CascadeMux I__9100 (
            .O(N__37474),
            .I(N__37459));
    InMux I__9099 (
            .O(N__37471),
            .I(N__37456));
    LocalMux I__9098 (
            .O(N__37468),
            .I(N__37453));
    InMux I__9097 (
            .O(N__37467),
            .I(N__37450));
    InMux I__9096 (
            .O(N__37466),
            .I(N__37445));
    InMux I__9095 (
            .O(N__37463),
            .I(N__37445));
    CascadeMux I__9094 (
            .O(N__37462),
            .I(N__37442));
    InMux I__9093 (
            .O(N__37459),
            .I(N__37438));
    LocalMux I__9092 (
            .O(N__37456),
            .I(N__37435));
    Span4Mux_v I__9091 (
            .O(N__37453),
            .I(N__37428));
    LocalMux I__9090 (
            .O(N__37450),
            .I(N__37428));
    LocalMux I__9089 (
            .O(N__37445),
            .I(N__37428));
    InMux I__9088 (
            .O(N__37442),
            .I(N__37425));
    CascadeMux I__9087 (
            .O(N__37441),
            .I(N__37422));
    LocalMux I__9086 (
            .O(N__37438),
            .I(N__37418));
    Span4Mux_v I__9085 (
            .O(N__37435),
            .I(N__37415));
    Span4Mux_v I__9084 (
            .O(N__37428),
            .I(N__37412));
    LocalMux I__9083 (
            .O(N__37425),
            .I(N__37409));
    InMux I__9082 (
            .O(N__37422),
            .I(N__37406));
    InMux I__9081 (
            .O(N__37421),
            .I(N__37403));
    Span4Mux_v I__9080 (
            .O(N__37418),
            .I(N__37400));
    Span4Mux_v I__9079 (
            .O(N__37415),
            .I(N__37391));
    Span4Mux_h I__9078 (
            .O(N__37412),
            .I(N__37391));
    Span4Mux_v I__9077 (
            .O(N__37409),
            .I(N__37391));
    LocalMux I__9076 (
            .O(N__37406),
            .I(N__37391));
    LocalMux I__9075 (
            .O(N__37403),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__9074 (
            .O(N__37400),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__9073 (
            .O(N__37391),
            .I(M_this_spr_address_qZ0Z_13));
    InMux I__9072 (
            .O(N__37384),
            .I(N__37380));
    CascadeMux I__9071 (
            .O(N__37383),
            .I(N__37376));
    LocalMux I__9070 (
            .O(N__37380),
            .I(N__37370));
    InMux I__9069 (
            .O(N__37379),
            .I(N__37367));
    InMux I__9068 (
            .O(N__37376),
            .I(N__37362));
    InMux I__9067 (
            .O(N__37375),
            .I(N__37362));
    InMux I__9066 (
            .O(N__37374),
            .I(N__37359));
    InMux I__9065 (
            .O(N__37373),
            .I(N__37355));
    Span4Mux_v I__9064 (
            .O(N__37370),
            .I(N__37348));
    LocalMux I__9063 (
            .O(N__37367),
            .I(N__37348));
    LocalMux I__9062 (
            .O(N__37362),
            .I(N__37348));
    LocalMux I__9061 (
            .O(N__37359),
            .I(N__37345));
    InMux I__9060 (
            .O(N__37358),
            .I(N__37342));
    LocalMux I__9059 (
            .O(N__37355),
            .I(N__37337));
    Span4Mux_v I__9058 (
            .O(N__37348),
            .I(N__37334));
    Span4Mux_v I__9057 (
            .O(N__37345),
            .I(N__37329));
    LocalMux I__9056 (
            .O(N__37342),
            .I(N__37329));
    InMux I__9055 (
            .O(N__37341),
            .I(N__37326));
    InMux I__9054 (
            .O(N__37340),
            .I(N__37323));
    Span4Mux_v I__9053 (
            .O(N__37337),
            .I(N__37320));
    Span4Mux_h I__9052 (
            .O(N__37334),
            .I(N__37313));
    Span4Mux_v I__9051 (
            .O(N__37329),
            .I(N__37313));
    LocalMux I__9050 (
            .O(N__37326),
            .I(N__37313));
    LocalMux I__9049 (
            .O(N__37323),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__9048 (
            .O(N__37320),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__9047 (
            .O(N__37313),
            .I(M_this_spr_address_qZ0Z_12));
    CascadeMux I__9046 (
            .O(N__37306),
            .I(N__37297));
    CascadeMux I__9045 (
            .O(N__37305),
            .I(N__37294));
    InMux I__9044 (
            .O(N__37304),
            .I(N__37291));
    InMux I__9043 (
            .O(N__37303),
            .I(N__37288));
    InMux I__9042 (
            .O(N__37302),
            .I(N__37283));
    InMux I__9041 (
            .O(N__37301),
            .I(N__37283));
    InMux I__9040 (
            .O(N__37300),
            .I(N__37280));
    InMux I__9039 (
            .O(N__37297),
            .I(N__37277));
    InMux I__9038 (
            .O(N__37294),
            .I(N__37274));
    LocalMux I__9037 (
            .O(N__37291),
            .I(N__37270));
    LocalMux I__9036 (
            .O(N__37288),
            .I(N__37267));
    LocalMux I__9035 (
            .O(N__37283),
            .I(N__37264));
    LocalMux I__9034 (
            .O(N__37280),
            .I(N__37261));
    LocalMux I__9033 (
            .O(N__37277),
            .I(N__37255));
    LocalMux I__9032 (
            .O(N__37274),
            .I(N__37255));
    InMux I__9031 (
            .O(N__37273),
            .I(N__37252));
    Span4Mux_v I__9030 (
            .O(N__37270),
            .I(N__37249));
    Span4Mux_v I__9029 (
            .O(N__37267),
            .I(N__37244));
    Span4Mux_h I__9028 (
            .O(N__37264),
            .I(N__37244));
    Span4Mux_h I__9027 (
            .O(N__37261),
            .I(N__37241));
    InMux I__9026 (
            .O(N__37260),
            .I(N__37238));
    Span12Mux_v I__9025 (
            .O(N__37255),
            .I(N__37233));
    LocalMux I__9024 (
            .O(N__37252),
            .I(N__37233));
    Span4Mux_h I__9023 (
            .O(N__37249),
            .I(N__37230));
    Span4Mux_h I__9022 (
            .O(N__37244),
            .I(N__37225));
    Span4Mux_v I__9021 (
            .O(N__37241),
            .I(N__37225));
    LocalMux I__9020 (
            .O(N__37238),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv12 I__9019 (
            .O(N__37233),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__9018 (
            .O(N__37230),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__9017 (
            .O(N__37225),
            .I(M_this_spr_address_qZ0Z_11));
    CEMux I__9016 (
            .O(N__37216),
            .I(N__37213));
    LocalMux I__9015 (
            .O(N__37213),
            .I(N__37209));
    CEMux I__9014 (
            .O(N__37212),
            .I(N__37206));
    Odrv4 I__9013 (
            .O(N__37209),
            .I(\this_spr_ram.mem_WE_12 ));
    LocalMux I__9012 (
            .O(N__37206),
            .I(\this_spr_ram.mem_WE_12 ));
    InMux I__9011 (
            .O(N__37201),
            .I(N__37198));
    LocalMux I__9010 (
            .O(N__37198),
            .I(N__37195));
    Span4Mux_v I__9009 (
            .O(N__37195),
            .I(N__37190));
    InMux I__9008 (
            .O(N__37194),
            .I(N__37187));
    InMux I__9007 (
            .O(N__37193),
            .I(N__37184));
    Sp12to4 I__9006 (
            .O(N__37190),
            .I(N__37178));
    LocalMux I__9005 (
            .O(N__37187),
            .I(N__37178));
    LocalMux I__9004 (
            .O(N__37184),
            .I(N__37175));
    InMux I__9003 (
            .O(N__37183),
            .I(N__37172));
    Odrv12 I__9002 (
            .O(N__37178),
            .I(\this_ppu.N_545 ));
    Odrv4 I__9001 (
            .O(N__37175),
            .I(\this_ppu.N_545 ));
    LocalMux I__9000 (
            .O(N__37172),
            .I(\this_ppu.N_545 ));
    InMux I__8999 (
            .O(N__37165),
            .I(N__37162));
    LocalMux I__8998 (
            .O(N__37162),
            .I(N__37158));
    InMux I__8997 (
            .O(N__37161),
            .I(N__37155));
    Span4Mux_h I__8996 (
            .O(N__37158),
            .I(N__37150));
    LocalMux I__8995 (
            .O(N__37155),
            .I(N__37147));
    InMux I__8994 (
            .O(N__37154),
            .I(N__37144));
    InMux I__8993 (
            .O(N__37153),
            .I(N__37141));
    Span4Mux_v I__8992 (
            .O(N__37150),
            .I(N__37135));
    Span4Mux_h I__8991 (
            .O(N__37147),
            .I(N__37135));
    LocalMux I__8990 (
            .O(N__37144),
            .I(N__37132));
    LocalMux I__8989 (
            .O(N__37141),
            .I(N__37129));
    InMux I__8988 (
            .O(N__37140),
            .I(N__37126));
    Span4Mux_v I__8987 (
            .O(N__37135),
            .I(N__37120));
    Span4Mux_h I__8986 (
            .O(N__37132),
            .I(N__37120));
    Span4Mux_s2_v I__8985 (
            .O(N__37129),
            .I(N__37115));
    LocalMux I__8984 (
            .O(N__37126),
            .I(N__37115));
    InMux I__8983 (
            .O(N__37125),
            .I(N__37112));
    Sp12to4 I__8982 (
            .O(N__37120),
            .I(N__37108));
    Span4Mux_v I__8981 (
            .O(N__37115),
            .I(N__37103));
    LocalMux I__8980 (
            .O(N__37112),
            .I(N__37103));
    InMux I__8979 (
            .O(N__37111),
            .I(N__37100));
    Span12Mux_h I__8978 (
            .O(N__37108),
            .I(N__37096));
    Span4Mux_v I__8977 (
            .O(N__37103),
            .I(N__37093));
    LocalMux I__8976 (
            .O(N__37100),
            .I(N__37090));
    InMux I__8975 (
            .O(N__37099),
            .I(N__37087));
    Odrv12 I__8974 (
            .O(N__37096),
            .I(M_this_spr_ram_write_data_3));
    Odrv4 I__8973 (
            .O(N__37093),
            .I(M_this_spr_ram_write_data_3));
    Odrv4 I__8972 (
            .O(N__37090),
            .I(M_this_spr_ram_write_data_3));
    LocalMux I__8971 (
            .O(N__37087),
            .I(M_this_spr_ram_write_data_3));
    InMux I__8970 (
            .O(N__37078),
            .I(N__37071));
    CascadeMux I__8969 (
            .O(N__37077),
            .I(N__37068));
    CascadeMux I__8968 (
            .O(N__37076),
            .I(N__37065));
    InMux I__8967 (
            .O(N__37075),
            .I(N__37058));
    InMux I__8966 (
            .O(N__37074),
            .I(N__37058));
    LocalMux I__8965 (
            .O(N__37071),
            .I(N__37055));
    InMux I__8964 (
            .O(N__37068),
            .I(N__37052));
    InMux I__8963 (
            .O(N__37065),
            .I(N__37049));
    InMux I__8962 (
            .O(N__37064),
            .I(N__37046));
    InMux I__8961 (
            .O(N__37063),
            .I(N__37043));
    LocalMux I__8960 (
            .O(N__37058),
            .I(N__37040));
    Span4Mux_v I__8959 (
            .O(N__37055),
            .I(N__37033));
    LocalMux I__8958 (
            .O(N__37052),
            .I(N__37033));
    LocalMux I__8957 (
            .O(N__37049),
            .I(N__37033));
    LocalMux I__8956 (
            .O(N__37046),
            .I(N__37030));
    LocalMux I__8955 (
            .O(N__37043),
            .I(N__37027));
    Span4Mux_v I__8954 (
            .O(N__37040),
            .I(N__37024));
    Span4Mux_h I__8953 (
            .O(N__37033),
            .I(N__37021));
    Span4Mux_v I__8952 (
            .O(N__37030),
            .I(N__37018));
    Span4Mux_v I__8951 (
            .O(N__37027),
            .I(N__37015));
    Span4Mux_v I__8950 (
            .O(N__37024),
            .I(N__37012));
    Sp12to4 I__8949 (
            .O(N__37021),
            .I(N__37009));
    Span4Mux_h I__8948 (
            .O(N__37018),
            .I(N__37004));
    Span4Mux_v I__8947 (
            .O(N__37015),
            .I(N__37004));
    Sp12to4 I__8946 (
            .O(N__37012),
            .I(N__37001));
    Span12Mux_v I__8945 (
            .O(N__37009),
            .I(N__36998));
    Span4Mux_h I__8944 (
            .O(N__37004),
            .I(N__36995));
    Odrv12 I__8943 (
            .O(N__37001),
            .I(port_address_in_4));
    Odrv12 I__8942 (
            .O(N__36998),
            .I(port_address_in_4));
    Odrv4 I__8941 (
            .O(N__36995),
            .I(port_address_in_4));
    InMux I__8940 (
            .O(N__36988),
            .I(N__36982));
    InMux I__8939 (
            .O(N__36987),
            .I(N__36977));
    InMux I__8938 (
            .O(N__36986),
            .I(N__36977));
    InMux I__8937 (
            .O(N__36985),
            .I(N__36974));
    LocalMux I__8936 (
            .O(N__36982),
            .I(N__36968));
    LocalMux I__8935 (
            .O(N__36977),
            .I(N__36968));
    LocalMux I__8934 (
            .O(N__36974),
            .I(N__36963));
    InMux I__8933 (
            .O(N__36973),
            .I(N__36960));
    Span4Mux_v I__8932 (
            .O(N__36968),
            .I(N__36957));
    InMux I__8931 (
            .O(N__36967),
            .I(N__36954));
    InMux I__8930 (
            .O(N__36966),
            .I(N__36951));
    Span4Mux_v I__8929 (
            .O(N__36963),
            .I(N__36946));
    LocalMux I__8928 (
            .O(N__36960),
            .I(N__36946));
    Sp12to4 I__8927 (
            .O(N__36957),
            .I(N__36939));
    LocalMux I__8926 (
            .O(N__36954),
            .I(N__36939));
    LocalMux I__8925 (
            .O(N__36951),
            .I(N__36939));
    Span4Mux_v I__8924 (
            .O(N__36946),
            .I(N__36936));
    Span12Mux_h I__8923 (
            .O(N__36939),
            .I(N__36933));
    Span4Mux_h I__8922 (
            .O(N__36936),
            .I(N__36930));
    Span12Mux_v I__8921 (
            .O(N__36933),
            .I(N__36927));
    Sp12to4 I__8920 (
            .O(N__36930),
            .I(N__36924));
    Odrv12 I__8919 (
            .O(N__36927),
            .I(port_address_in_0));
    Odrv12 I__8918 (
            .O(N__36924),
            .I(port_address_in_0));
    CascadeMux I__8917 (
            .O(N__36919),
            .I(N__36916));
    InMux I__8916 (
            .O(N__36916),
            .I(N__36913));
    LocalMux I__8915 (
            .O(N__36913),
            .I(\this_ppu.N_610 ));
    InMux I__8914 (
            .O(N__36910),
            .I(N__36907));
    LocalMux I__8913 (
            .O(N__36907),
            .I(M_this_state_d_0_sqmuxa_2));
    IoInMux I__8912 (
            .O(N__36904),
            .I(N__36901));
    LocalMux I__8911 (
            .O(N__36901),
            .I(N__36898));
    IoSpan4Mux I__8910 (
            .O(N__36898),
            .I(N__36895));
    Span4Mux_s0_h I__8909 (
            .O(N__36895),
            .I(N__36890));
    CascadeMux I__8908 (
            .O(N__36894),
            .I(N__36887));
    CascadeMux I__8907 (
            .O(N__36893),
            .I(N__36882));
    Sp12to4 I__8906 (
            .O(N__36890),
            .I(N__36879));
    InMux I__8905 (
            .O(N__36887),
            .I(N__36876));
    InMux I__8904 (
            .O(N__36886),
            .I(N__36872));
    InMux I__8903 (
            .O(N__36885),
            .I(N__36867));
    InMux I__8902 (
            .O(N__36882),
            .I(N__36867));
    Span12Mux_v I__8901 (
            .O(N__36879),
            .I(N__36864));
    LocalMux I__8900 (
            .O(N__36876),
            .I(N__36861));
    InMux I__8899 (
            .O(N__36875),
            .I(N__36858));
    LocalMux I__8898 (
            .O(N__36872),
            .I(N__36853));
    LocalMux I__8897 (
            .O(N__36867),
            .I(N__36853));
    Odrv12 I__8896 (
            .O(N__36864),
            .I(led_c_1));
    Odrv4 I__8895 (
            .O(N__36861),
            .I(led_c_1));
    LocalMux I__8894 (
            .O(N__36858),
            .I(led_c_1));
    Odrv4 I__8893 (
            .O(N__36853),
            .I(led_c_1));
    InMux I__8892 (
            .O(N__36844),
            .I(N__36840));
    InMux I__8891 (
            .O(N__36843),
            .I(N__36837));
    LocalMux I__8890 (
            .O(N__36840),
            .I(N_608));
    LocalMux I__8889 (
            .O(N__36837),
            .I(N_608));
    InMux I__8888 (
            .O(N__36832),
            .I(N__36826));
    InMux I__8887 (
            .O(N__36831),
            .I(N__36821));
    InMux I__8886 (
            .O(N__36830),
            .I(N__36821));
    InMux I__8885 (
            .O(N__36829),
            .I(N__36818));
    LocalMux I__8884 (
            .O(N__36826),
            .I(M_this_substate_qZ0));
    LocalMux I__8883 (
            .O(N__36821),
            .I(M_this_substate_qZ0));
    LocalMux I__8882 (
            .O(N__36818),
            .I(M_this_substate_qZ0));
    CascadeMux I__8881 (
            .O(N__36811),
            .I(N__36807));
    InMux I__8880 (
            .O(N__36810),
            .I(N__36803));
    InMux I__8879 (
            .O(N__36807),
            .I(N__36800));
    CascadeMux I__8878 (
            .O(N__36806),
            .I(N__36793));
    LocalMux I__8877 (
            .O(N__36803),
            .I(N__36790));
    LocalMux I__8876 (
            .O(N__36800),
            .I(N__36787));
    InMux I__8875 (
            .O(N__36799),
            .I(N__36784));
    CascadeMux I__8874 (
            .O(N__36798),
            .I(N__36781));
    CascadeMux I__8873 (
            .O(N__36797),
            .I(N__36778));
    InMux I__8872 (
            .O(N__36796),
            .I(N__36770));
    InMux I__8871 (
            .O(N__36793),
            .I(N__36770));
    Span4Mux_v I__8870 (
            .O(N__36790),
            .I(N__36767));
    Span12Mux_v I__8869 (
            .O(N__36787),
            .I(N__36762));
    LocalMux I__8868 (
            .O(N__36784),
            .I(N__36762));
    InMux I__8867 (
            .O(N__36781),
            .I(N__36757));
    InMux I__8866 (
            .O(N__36778),
            .I(N__36757));
    InMux I__8865 (
            .O(N__36777),
            .I(N__36750));
    InMux I__8864 (
            .O(N__36776),
            .I(N__36750));
    InMux I__8863 (
            .O(N__36775),
            .I(N__36750));
    LocalMux I__8862 (
            .O(N__36770),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8861 (
            .O(N__36767),
            .I(M_this_state_qZ0Z_13));
    Odrv12 I__8860 (
            .O(N__36762),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__8859 (
            .O(N__36757),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__8858 (
            .O(N__36750),
            .I(M_this_state_qZ0Z_13));
    InMux I__8857 (
            .O(N__36739),
            .I(N__36735));
    InMux I__8856 (
            .O(N__36738),
            .I(N__36732));
    LocalMux I__8855 (
            .O(N__36735),
            .I(N__36728));
    LocalMux I__8854 (
            .O(N__36732),
            .I(N__36723));
    InMux I__8853 (
            .O(N__36731),
            .I(N__36718));
    Span4Mux_h I__8852 (
            .O(N__36728),
            .I(N__36715));
    InMux I__8851 (
            .O(N__36727),
            .I(N__36710));
    InMux I__8850 (
            .O(N__36726),
            .I(N__36710));
    Span4Mux_v I__8849 (
            .O(N__36723),
            .I(N__36707));
    InMux I__8848 (
            .O(N__36722),
            .I(N__36704));
    InMux I__8847 (
            .O(N__36721),
            .I(N__36701));
    LocalMux I__8846 (
            .O(N__36718),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__8845 (
            .O(N__36715),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__8844 (
            .O(N__36710),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__8843 (
            .O(N__36707),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__8842 (
            .O(N__36704),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__8841 (
            .O(N__36701),
            .I(M_this_state_qZ0Z_11));
    InMux I__8840 (
            .O(N__36688),
            .I(N__36684));
    CascadeMux I__8839 (
            .O(N__36687),
            .I(N__36680));
    LocalMux I__8838 (
            .O(N__36684),
            .I(N__36674));
    InMux I__8837 (
            .O(N__36683),
            .I(N__36671));
    InMux I__8836 (
            .O(N__36680),
            .I(N__36664));
    InMux I__8835 (
            .O(N__36679),
            .I(N__36661));
    InMux I__8834 (
            .O(N__36678),
            .I(N__36658));
    InMux I__8833 (
            .O(N__36677),
            .I(N__36653));
    Span4Mux_h I__8832 (
            .O(N__36674),
            .I(N__36648));
    LocalMux I__8831 (
            .O(N__36671),
            .I(N__36648));
    InMux I__8830 (
            .O(N__36670),
            .I(N__36643));
    InMux I__8829 (
            .O(N__36669),
            .I(N__36643));
    InMux I__8828 (
            .O(N__36668),
            .I(N__36638));
    InMux I__8827 (
            .O(N__36667),
            .I(N__36638));
    LocalMux I__8826 (
            .O(N__36664),
            .I(N__36635));
    LocalMux I__8825 (
            .O(N__36661),
            .I(N__36632));
    LocalMux I__8824 (
            .O(N__36658),
            .I(N__36629));
    InMux I__8823 (
            .O(N__36657),
            .I(N__36626));
    InMux I__8822 (
            .O(N__36656),
            .I(N__36623));
    LocalMux I__8821 (
            .O(N__36653),
            .I(N__36618));
    Span4Mux_h I__8820 (
            .O(N__36648),
            .I(N__36618));
    LocalMux I__8819 (
            .O(N__36643),
            .I(N__36613));
    LocalMux I__8818 (
            .O(N__36638),
            .I(N__36613));
    Span12Mux_h I__8817 (
            .O(N__36635),
            .I(N__36610));
    Odrv12 I__8816 (
            .O(N__36632),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__8815 (
            .O(N__36629),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__8814 (
            .O(N__36626),
            .I(M_this_state_qZ0Z_9));
    LocalMux I__8813 (
            .O(N__36623),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__8812 (
            .O(N__36618),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__8811 (
            .O(N__36613),
            .I(M_this_state_qZ0Z_9));
    Odrv12 I__8810 (
            .O(N__36610),
            .I(M_this_state_qZ0Z_9));
    InMux I__8809 (
            .O(N__36595),
            .I(N__36592));
    LocalMux I__8808 (
            .O(N__36592),
            .I(N__36589));
    Odrv4 I__8807 (
            .O(N__36589),
            .I(\this_ppu.oam_cache.mem_10 ));
    CascadeMux I__8806 (
            .O(N__36586),
            .I(N__36583));
    InMux I__8805 (
            .O(N__36583),
            .I(N__36578));
    InMux I__8804 (
            .O(N__36582),
            .I(N__36575));
    InMux I__8803 (
            .O(N__36581),
            .I(N__36572));
    LocalMux I__8802 (
            .O(N__36578),
            .I(N__36569));
    LocalMux I__8801 (
            .O(N__36575),
            .I(N__36563));
    LocalMux I__8800 (
            .O(N__36572),
            .I(N__36563));
    Span4Mux_h I__8799 (
            .O(N__36569),
            .I(N__36557));
    InMux I__8798 (
            .O(N__36568),
            .I(N__36554));
    Span4Mux_h I__8797 (
            .O(N__36563),
            .I(N__36551));
    InMux I__8796 (
            .O(N__36562),
            .I(N__36544));
    InMux I__8795 (
            .O(N__36561),
            .I(N__36544));
    InMux I__8794 (
            .O(N__36560),
            .I(N__36544));
    Odrv4 I__8793 (
            .O(N__36557),
            .I(\this_ppu.un1_M_hoffset_q_5 ));
    LocalMux I__8792 (
            .O(N__36554),
            .I(\this_ppu.un1_M_hoffset_q_5 ));
    Odrv4 I__8791 (
            .O(N__36551),
            .I(\this_ppu.un1_M_hoffset_q_5 ));
    LocalMux I__8790 (
            .O(N__36544),
            .I(\this_ppu.un1_M_hoffset_q_5 ));
    InMux I__8789 (
            .O(N__36535),
            .I(N__36532));
    LocalMux I__8788 (
            .O(N__36532),
            .I(N__36529));
    Span4Mux_v I__8787 (
            .O(N__36529),
            .I(N__36526));
    Odrv4 I__8786 (
            .O(N__36526),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_18 ));
    InMux I__8785 (
            .O(N__36523),
            .I(N__36520));
    LocalMux I__8784 (
            .O(N__36520),
            .I(N__36515));
    InMux I__8783 (
            .O(N__36519),
            .I(N__36512));
    CascadeMux I__8782 (
            .O(N__36518),
            .I(N__36509));
    Span4Mux_h I__8781 (
            .O(N__36515),
            .I(N__36505));
    LocalMux I__8780 (
            .O(N__36512),
            .I(N__36502));
    InMux I__8779 (
            .O(N__36509),
            .I(N__36499));
    InMux I__8778 (
            .O(N__36508),
            .I(N__36496));
    Odrv4 I__8777 (
            .O(N__36505),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__8776 (
            .O(N__36502),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__8775 (
            .O(N__36499),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__8774 (
            .O(N__36496),
            .I(M_this_state_qZ0Z_1));
    InMux I__8773 (
            .O(N__36487),
            .I(N__36482));
    InMux I__8772 (
            .O(N__36486),
            .I(N__36479));
    CascadeMux I__8771 (
            .O(N__36485),
            .I(N__36473));
    LocalMux I__8770 (
            .O(N__36482),
            .I(N__36469));
    LocalMux I__8769 (
            .O(N__36479),
            .I(N__36466));
    InMux I__8768 (
            .O(N__36478),
            .I(N__36463));
    InMux I__8767 (
            .O(N__36477),
            .I(N__36459));
    InMux I__8766 (
            .O(N__36476),
            .I(N__36453));
    InMux I__8765 (
            .O(N__36473),
            .I(N__36453));
    InMux I__8764 (
            .O(N__36472),
            .I(N__36450));
    Span4Mux_h I__8763 (
            .O(N__36469),
            .I(N__36445));
    Span4Mux_v I__8762 (
            .O(N__36466),
            .I(N__36445));
    LocalMux I__8761 (
            .O(N__36463),
            .I(N__36442));
    InMux I__8760 (
            .O(N__36462),
            .I(N__36439));
    LocalMux I__8759 (
            .O(N__36459),
            .I(N__36436));
    InMux I__8758 (
            .O(N__36458),
            .I(N__36433));
    LocalMux I__8757 (
            .O(N__36453),
            .I(N__36430));
    LocalMux I__8756 (
            .O(N__36450),
            .I(N__36426));
    Span4Mux_v I__8755 (
            .O(N__36445),
            .I(N__36423));
    Span4Mux_v I__8754 (
            .O(N__36442),
            .I(N__36420));
    LocalMux I__8753 (
            .O(N__36439),
            .I(N__36415));
    Span4Mux_h I__8752 (
            .O(N__36436),
            .I(N__36415));
    LocalMux I__8751 (
            .O(N__36433),
            .I(N__36412));
    Span4Mux_v I__8750 (
            .O(N__36430),
            .I(N__36409));
    InMux I__8749 (
            .O(N__36429),
            .I(N__36406));
    Span12Mux_s10_v I__8748 (
            .O(N__36426),
            .I(N__36403));
    Sp12to4 I__8747 (
            .O(N__36423),
            .I(N__36400));
    Sp12to4 I__8746 (
            .O(N__36420),
            .I(N__36397));
    Span4Mux_v I__8745 (
            .O(N__36415),
            .I(N__36394));
    Span4Mux_h I__8744 (
            .O(N__36412),
            .I(N__36391));
    Span4Mux_v I__8743 (
            .O(N__36409),
            .I(N__36388));
    LocalMux I__8742 (
            .O(N__36406),
            .I(N__36385));
    Span12Mux_v I__8741 (
            .O(N__36403),
            .I(N__36382));
    Span12Mux_h I__8740 (
            .O(N__36400),
            .I(N__36379));
    Span12Mux_h I__8739 (
            .O(N__36397),
            .I(N__36372));
    Sp12to4 I__8738 (
            .O(N__36394),
            .I(N__36372));
    Sp12to4 I__8737 (
            .O(N__36391),
            .I(N__36372));
    Span4Mux_v I__8736 (
            .O(N__36388),
            .I(N__36367));
    Span4Mux_v I__8735 (
            .O(N__36385),
            .I(N__36367));
    Span12Mux_h I__8734 (
            .O(N__36382),
            .I(N__36362));
    Span12Mux_v I__8733 (
            .O(N__36379),
            .I(N__36362));
    Span12Mux_v I__8732 (
            .O(N__36372),
            .I(N__36359));
    Span4Mux_h I__8731 (
            .O(N__36367),
            .I(N__36356));
    Odrv12 I__8730 (
            .O(N__36362),
            .I(port_data_c_7));
    Odrv12 I__8729 (
            .O(N__36359),
            .I(port_data_c_7));
    Odrv4 I__8728 (
            .O(N__36356),
            .I(port_data_c_7));
    InMux I__8727 (
            .O(N__36349),
            .I(N__36346));
    LocalMux I__8726 (
            .O(N__36346),
            .I(N__36343));
    Odrv4 I__8725 (
            .O(N__36343),
            .I(N_440));
    InMux I__8724 (
            .O(N__36340),
            .I(N__36337));
    LocalMux I__8723 (
            .O(N__36337),
            .I(N__36334));
    Odrv4 I__8722 (
            .O(N__36334),
            .I(N_437));
    InMux I__8721 (
            .O(N__36331),
            .I(N__36328));
    LocalMux I__8720 (
            .O(N__36328),
            .I(N__36325));
    Odrv4 I__8719 (
            .O(N__36325),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__8718 (
            .O(N__36322),
            .I(N__36319));
    LocalMux I__8717 (
            .O(N__36319),
            .I(N__36316));
    Odrv12 I__8716 (
            .O(N__36316),
            .I(M_this_oam_ram_write_data_22));
    InMux I__8715 (
            .O(N__36313),
            .I(N__36310));
    LocalMux I__8714 (
            .O(N__36310),
            .I(N__36304));
    InMux I__8713 (
            .O(N__36309),
            .I(N__36301));
    CascadeMux I__8712 (
            .O(N__36308),
            .I(N__36298));
    InMux I__8711 (
            .O(N__36307),
            .I(N__36295));
    Span4Mux_v I__8710 (
            .O(N__36304),
            .I(N__36288));
    LocalMux I__8709 (
            .O(N__36301),
            .I(N__36288));
    InMux I__8708 (
            .O(N__36298),
            .I(N__36285));
    LocalMux I__8707 (
            .O(N__36295),
            .I(N__36282));
    CascadeMux I__8706 (
            .O(N__36294),
            .I(N__36279));
    InMux I__8705 (
            .O(N__36293),
            .I(N__36275));
    Span4Mux_v I__8704 (
            .O(N__36288),
            .I(N__36270));
    LocalMux I__8703 (
            .O(N__36285),
            .I(N__36270));
    Span4Mux_v I__8702 (
            .O(N__36282),
            .I(N__36266));
    InMux I__8701 (
            .O(N__36279),
            .I(N__36263));
    InMux I__8700 (
            .O(N__36278),
            .I(N__36259));
    LocalMux I__8699 (
            .O(N__36275),
            .I(N__36256));
    Span4Mux_v I__8698 (
            .O(N__36270),
            .I(N__36253));
    InMux I__8697 (
            .O(N__36269),
            .I(N__36250));
    Span4Mux_v I__8696 (
            .O(N__36266),
            .I(N__36247));
    LocalMux I__8695 (
            .O(N__36263),
            .I(N__36244));
    InMux I__8694 (
            .O(N__36262),
            .I(N__36241));
    LocalMux I__8693 (
            .O(N__36259),
            .I(N__36238));
    Sp12to4 I__8692 (
            .O(N__36256),
            .I(N__36235));
    Span4Mux_h I__8691 (
            .O(N__36253),
            .I(N__36230));
    LocalMux I__8690 (
            .O(N__36250),
            .I(N__36230));
    Sp12to4 I__8689 (
            .O(N__36247),
            .I(N__36227));
    Span4Mux_v I__8688 (
            .O(N__36244),
            .I(N__36224));
    LocalMux I__8687 (
            .O(N__36241),
            .I(N__36221));
    Span12Mux_h I__8686 (
            .O(N__36238),
            .I(N__36214));
    Span12Mux_s9_v I__8685 (
            .O(N__36235),
            .I(N__36214));
    Sp12to4 I__8684 (
            .O(N__36230),
            .I(N__36214));
    Span12Mux_h I__8683 (
            .O(N__36227),
            .I(N__36211));
    Sp12to4 I__8682 (
            .O(N__36224),
            .I(N__36208));
    Span12Mux_h I__8681 (
            .O(N__36221),
            .I(N__36205));
    Span12Mux_v I__8680 (
            .O(N__36214),
            .I(N__36202));
    Span12Mux_v I__8679 (
            .O(N__36211),
            .I(N__36199));
    Span12Mux_h I__8678 (
            .O(N__36208),
            .I(N__36196));
    Span12Mux_v I__8677 (
            .O(N__36205),
            .I(N__36191));
    Span12Mux_h I__8676 (
            .O(N__36202),
            .I(N__36191));
    Odrv12 I__8675 (
            .O(N__36199),
            .I(port_data_c_6));
    Odrv12 I__8674 (
            .O(N__36196),
            .I(port_data_c_6));
    Odrv12 I__8673 (
            .O(N__36191),
            .I(port_data_c_6));
    InMux I__8672 (
            .O(N__36184),
            .I(N__36181));
    LocalMux I__8671 (
            .O(N__36181),
            .I(N__36178));
    Span4Mux_h I__8670 (
            .O(N__36178),
            .I(N__36175));
    Odrv4 I__8669 (
            .O(N__36175),
            .I(N_439));
    CEMux I__8668 (
            .O(N__36172),
            .I(N__36169));
    LocalMux I__8667 (
            .O(N__36169),
            .I(N__36165));
    CEMux I__8666 (
            .O(N__36168),
            .I(N__36162));
    Odrv4 I__8665 (
            .O(N__36165),
            .I(\this_spr_ram.mem_WE_2 ));
    LocalMux I__8664 (
            .O(N__36162),
            .I(\this_spr_ram.mem_WE_2 ));
    CEMux I__8663 (
            .O(N__36157),
            .I(N__36153));
    CEMux I__8662 (
            .O(N__36156),
            .I(N__36150));
    LocalMux I__8661 (
            .O(N__36153),
            .I(\this_spr_ram.mem_WE_4 ));
    LocalMux I__8660 (
            .O(N__36150),
            .I(\this_spr_ram.mem_WE_4 ));
    InMux I__8659 (
            .O(N__36145),
            .I(N__36142));
    LocalMux I__8658 (
            .O(N__36142),
            .I(\this_spr_ram.mem_out_bus5_1 ));
    InMux I__8657 (
            .O(N__36139),
            .I(N__36136));
    LocalMux I__8656 (
            .O(N__36136),
            .I(N__36133));
    Span4Mux_h I__8655 (
            .O(N__36133),
            .I(N__36130));
    Odrv4 I__8654 (
            .O(N__36130),
            .I(\this_spr_ram.mem_out_bus1_1 ));
    InMux I__8653 (
            .O(N__36127),
            .I(N__36124));
    LocalMux I__8652 (
            .O(N__36124),
            .I(N__36121));
    Span12Mux_s10_v I__8651 (
            .O(N__36121),
            .I(N__36118));
    Odrv12 I__8650 (
            .O(N__36118),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ));
    CEMux I__8649 (
            .O(N__36115),
            .I(N__36111));
    CEMux I__8648 (
            .O(N__36114),
            .I(N__36108));
    LocalMux I__8647 (
            .O(N__36111),
            .I(N__36105));
    LocalMux I__8646 (
            .O(N__36108),
            .I(N__36102));
    Span4Mux_v I__8645 (
            .O(N__36105),
            .I(N__36099));
    Span4Mux_h I__8644 (
            .O(N__36102),
            .I(N__36096));
    Span4Mux_v I__8643 (
            .O(N__36099),
            .I(N__36093));
    Span4Mux_v I__8642 (
            .O(N__36096),
            .I(N__36090));
    Odrv4 I__8641 (
            .O(N__36093),
            .I(\this_spr_ram.mem_WE_14 ));
    Odrv4 I__8640 (
            .O(N__36090),
            .I(\this_spr_ram.mem_WE_14 ));
    InMux I__8639 (
            .O(N__36085),
            .I(N__36082));
    LocalMux I__8638 (
            .O(N__36082),
            .I(N__36079));
    Span4Mux_v I__8637 (
            .O(N__36079),
            .I(N__36076));
    Odrv4 I__8636 (
            .O(N__36076),
            .I(M_this_oam_ram_write_data_7));
    InMux I__8635 (
            .O(N__36073),
            .I(N__36070));
    LocalMux I__8634 (
            .O(N__36070),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__8633 (
            .O(N__36067),
            .I(N__36064));
    LocalMux I__8632 (
            .O(N__36064),
            .I(N__36061));
    Span4Mux_h I__8631 (
            .O(N__36061),
            .I(N__36058));
    Odrv4 I__8630 (
            .O(N__36058),
            .I(M_this_oam_ram_write_data_3));
    InMux I__8629 (
            .O(N__36055),
            .I(N__36052));
    LocalMux I__8628 (
            .O(N__36052),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__8627 (
            .O(N__36049),
            .I(N__36046));
    LocalMux I__8626 (
            .O(N__36046),
            .I(N__36043));
    Span4Mux_h I__8625 (
            .O(N__36043),
            .I(N__36040));
    Odrv4 I__8624 (
            .O(N__36040),
            .I(M_this_oam_ram_write_data_4));
    InMux I__8623 (
            .O(N__36037),
            .I(N__36034));
    LocalMux I__8622 (
            .O(N__36034),
            .I(M_this_data_tmp_qZ0Z_4));
    CEMux I__8621 (
            .O(N__36031),
            .I(N__36025));
    CEMux I__8620 (
            .O(N__36030),
            .I(N__36022));
    CEMux I__8619 (
            .O(N__36029),
            .I(N__36019));
    CEMux I__8618 (
            .O(N__36028),
            .I(N__36016));
    LocalMux I__8617 (
            .O(N__36025),
            .I(N__36012));
    LocalMux I__8616 (
            .O(N__36022),
            .I(N__36009));
    LocalMux I__8615 (
            .O(N__36019),
            .I(N__36004));
    LocalMux I__8614 (
            .O(N__36016),
            .I(N__36004));
    CEMux I__8613 (
            .O(N__36015),
            .I(N__36001));
    Span4Mux_v I__8612 (
            .O(N__36012),
            .I(N__35998));
    Span4Mux_h I__8611 (
            .O(N__36009),
            .I(N__35995));
    Span4Mux_v I__8610 (
            .O(N__36004),
            .I(N__35990));
    LocalMux I__8609 (
            .O(N__36001),
            .I(N__35990));
    Span4Mux_h I__8608 (
            .O(N__35998),
            .I(N__35987));
    Span4Mux_h I__8607 (
            .O(N__35995),
            .I(N__35984));
    Span4Mux_h I__8606 (
            .O(N__35990),
            .I(N__35981));
    Odrv4 I__8605 (
            .O(N__35987),
            .I(N_1302_0));
    Odrv4 I__8604 (
            .O(N__35984),
            .I(N_1302_0));
    Odrv4 I__8603 (
            .O(N__35981),
            .I(N_1302_0));
    InMux I__8602 (
            .O(N__35974),
            .I(N__35971));
    LocalMux I__8601 (
            .O(N__35971),
            .I(N__35968));
    Odrv12 I__8600 (
            .O(N__35968),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__8599 (
            .O(N__35965),
            .I(N__35962));
    LocalMux I__8598 (
            .O(N__35962),
            .I(N__35959));
    Span4Mux_v I__8597 (
            .O(N__35959),
            .I(N__35956));
    Odrv4 I__8596 (
            .O(N__35956),
            .I(M_this_oam_ram_write_data_23));
    InMux I__8595 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__8594 (
            .O(N__35950),
            .I(N__35947));
    Span4Mux_v I__8593 (
            .O(N__35947),
            .I(N__35944));
    Odrv4 I__8592 (
            .O(N__35944),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_17 ));
    InMux I__8591 (
            .O(N__35941),
            .I(N__35938));
    LocalMux I__8590 (
            .O(N__35938),
            .I(N__35935));
    Odrv12 I__8589 (
            .O(N__35935),
            .I(\this_ppu.oam_cache.mem_11 ));
    InMux I__8588 (
            .O(N__35932),
            .I(N__35928));
    InMux I__8587 (
            .O(N__35931),
            .I(N__35925));
    LocalMux I__8586 (
            .O(N__35928),
            .I(N__35918));
    LocalMux I__8585 (
            .O(N__35925),
            .I(N__35918));
    CascadeMux I__8584 (
            .O(N__35924),
            .I(N__35915));
    CascadeMux I__8583 (
            .O(N__35923),
            .I(N__35912));
    Span4Mux_h I__8582 (
            .O(N__35918),
            .I(N__35909));
    InMux I__8581 (
            .O(N__35915),
            .I(N__35904));
    InMux I__8580 (
            .O(N__35912),
            .I(N__35904));
    Odrv4 I__8579 (
            .O(N__35909),
            .I(\this_ppu.un1_M_hoffset_q_6 ));
    LocalMux I__8578 (
            .O(N__35904),
            .I(\this_ppu.un1_M_hoffset_q_6 ));
    InMux I__8577 (
            .O(N__35899),
            .I(N__35894));
    InMux I__8576 (
            .O(N__35898),
            .I(N__35891));
    InMux I__8575 (
            .O(N__35897),
            .I(N__35888));
    LocalMux I__8574 (
            .O(N__35894),
            .I(N__35878));
    LocalMux I__8573 (
            .O(N__35891),
            .I(N__35878));
    LocalMux I__8572 (
            .O(N__35888),
            .I(N__35878));
    InMux I__8571 (
            .O(N__35887),
            .I(N__35875));
    InMux I__8570 (
            .O(N__35886),
            .I(N__35872));
    InMux I__8569 (
            .O(N__35885),
            .I(N__35869));
    Span4Mux_v I__8568 (
            .O(N__35878),
            .I(N__35864));
    LocalMux I__8567 (
            .O(N__35875),
            .I(N__35864));
    LocalMux I__8566 (
            .O(N__35872),
            .I(N__35861));
    LocalMux I__8565 (
            .O(N__35869),
            .I(N__35858));
    Span4Mux_h I__8564 (
            .O(N__35864),
            .I(N__35855));
    Odrv4 I__8563 (
            .O(N__35861),
            .I(\this_ppu.M_hoffset_qZ0Z_1 ));
    Odrv4 I__8562 (
            .O(N__35858),
            .I(\this_ppu.M_hoffset_qZ0Z_1 ));
    Odrv4 I__8561 (
            .O(N__35855),
            .I(\this_ppu.M_hoffset_qZ0Z_1 ));
    InMux I__8560 (
            .O(N__35848),
            .I(N__35843));
    InMux I__8559 (
            .O(N__35847),
            .I(N__35840));
    InMux I__8558 (
            .O(N__35846),
            .I(N__35837));
    LocalMux I__8557 (
            .O(N__35843),
            .I(N__35833));
    LocalMux I__8556 (
            .O(N__35840),
            .I(N__35827));
    LocalMux I__8555 (
            .O(N__35837),
            .I(N__35827));
    CascadeMux I__8554 (
            .O(N__35836),
            .I(N__35821));
    Span4Mux_h I__8553 (
            .O(N__35833),
            .I(N__35817));
    InMux I__8552 (
            .O(N__35832),
            .I(N__35814));
    Span4Mux_h I__8551 (
            .O(N__35827),
            .I(N__35811));
    InMux I__8550 (
            .O(N__35826),
            .I(N__35808));
    InMux I__8549 (
            .O(N__35825),
            .I(N__35805));
    InMux I__8548 (
            .O(N__35824),
            .I(N__35798));
    InMux I__8547 (
            .O(N__35821),
            .I(N__35798));
    InMux I__8546 (
            .O(N__35820),
            .I(N__35798));
    Odrv4 I__8545 (
            .O(N__35817),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    LocalMux I__8544 (
            .O(N__35814),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    Odrv4 I__8543 (
            .O(N__35811),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    LocalMux I__8542 (
            .O(N__35808),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    LocalMux I__8541 (
            .O(N__35805),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    LocalMux I__8540 (
            .O(N__35798),
            .I(\this_ppu.un1_M_hoffset_q_4 ));
    InMux I__8539 (
            .O(N__35785),
            .I(N__35778));
    InMux I__8538 (
            .O(N__35784),
            .I(N__35775));
    InMux I__8537 (
            .O(N__35783),
            .I(N__35772));
    InMux I__8536 (
            .O(N__35782),
            .I(N__35769));
    InMux I__8535 (
            .O(N__35781),
            .I(N__35766));
    LocalMux I__8534 (
            .O(N__35778),
            .I(N__35763));
    LocalMux I__8533 (
            .O(N__35775),
            .I(N__35754));
    LocalMux I__8532 (
            .O(N__35772),
            .I(N__35754));
    LocalMux I__8531 (
            .O(N__35769),
            .I(N__35754));
    LocalMux I__8530 (
            .O(N__35766),
            .I(N__35746));
    Span4Mux_h I__8529 (
            .O(N__35763),
            .I(N__35743));
    InMux I__8528 (
            .O(N__35762),
            .I(N__35740));
    InMux I__8527 (
            .O(N__35761),
            .I(N__35737));
    Span4Mux_v I__8526 (
            .O(N__35754),
            .I(N__35734));
    InMux I__8525 (
            .O(N__35753),
            .I(N__35731));
    InMux I__8524 (
            .O(N__35752),
            .I(N__35728));
    InMux I__8523 (
            .O(N__35751),
            .I(N__35721));
    InMux I__8522 (
            .O(N__35750),
            .I(N__35721));
    InMux I__8521 (
            .O(N__35749),
            .I(N__35721));
    Odrv12 I__8520 (
            .O(N__35746),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    Odrv4 I__8519 (
            .O(N__35743),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    LocalMux I__8518 (
            .O(N__35740),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    LocalMux I__8517 (
            .O(N__35737),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    Odrv4 I__8516 (
            .O(N__35734),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    LocalMux I__8515 (
            .O(N__35731),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    LocalMux I__8514 (
            .O(N__35728),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    LocalMux I__8513 (
            .O(N__35721),
            .I(\this_ppu.un1_M_hoffset_q_0 ));
    CascadeMux I__8512 (
            .O(N__35704),
            .I(N__35701));
    InMux I__8511 (
            .O(N__35701),
            .I(N__35698));
    LocalMux I__8510 (
            .O(N__35698),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0 ));
    InMux I__8509 (
            .O(N__35695),
            .I(N__35683));
    InMux I__8508 (
            .O(N__35694),
            .I(N__35683));
    InMux I__8507 (
            .O(N__35693),
            .I(N__35683));
    InMux I__8506 (
            .O(N__35692),
            .I(N__35683));
    LocalMux I__8505 (
            .O(N__35683),
            .I(\this_ppu.un1_oam_data_1_4_c5_0 ));
    CascadeMux I__8504 (
            .O(N__35680),
            .I(N__35676));
    InMux I__8503 (
            .O(N__35679),
            .I(N__35672));
    InMux I__8502 (
            .O(N__35676),
            .I(N__35666));
    InMux I__8501 (
            .O(N__35675),
            .I(N__35666));
    LocalMux I__8500 (
            .O(N__35672),
            .I(N__35663));
    InMux I__8499 (
            .O(N__35671),
            .I(N__35660));
    LocalMux I__8498 (
            .O(N__35666),
            .I(N__35657));
    Span4Mux_h I__8497 (
            .O(N__35663),
            .I(N__35654));
    LocalMux I__8496 (
            .O(N__35660),
            .I(N__35651));
    Span4Mux_h I__8495 (
            .O(N__35657),
            .I(N__35648));
    Span4Mux_v I__8494 (
            .O(N__35654),
            .I(N__35645));
    Span4Mux_h I__8493 (
            .O(N__35651),
            .I(N__35640));
    Span4Mux_v I__8492 (
            .O(N__35648),
            .I(N__35640));
    Odrv4 I__8491 (
            .O(N__35645),
            .I(M_this_oam_ram_read_data_23));
    Odrv4 I__8490 (
            .O(N__35640),
            .I(M_this_oam_ram_read_data_23));
    InMux I__8489 (
            .O(N__35635),
            .I(N__35632));
    LocalMux I__8488 (
            .O(N__35632),
            .I(N__35629));
    Span4Mux_h I__8487 (
            .O(N__35629),
            .I(N__35626));
    Odrv4 I__8486 (
            .O(N__35626),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_23 ));
    InMux I__8485 (
            .O(N__35623),
            .I(N__35620));
    LocalMux I__8484 (
            .O(N__35620),
            .I(N__35615));
    InMux I__8483 (
            .O(N__35619),
            .I(N__35612));
    CascadeMux I__8482 (
            .O(N__35618),
            .I(N__35609));
    Span4Mux_h I__8481 (
            .O(N__35615),
            .I(N__35603));
    LocalMux I__8480 (
            .O(N__35612),
            .I(N__35603));
    InMux I__8479 (
            .O(N__35609),
            .I(N__35599));
    InMux I__8478 (
            .O(N__35608),
            .I(N__35595));
    Span4Mux_h I__8477 (
            .O(N__35603),
            .I(N__35592));
    InMux I__8476 (
            .O(N__35602),
            .I(N__35589));
    LocalMux I__8475 (
            .O(N__35599),
            .I(N__35585));
    InMux I__8474 (
            .O(N__35598),
            .I(N__35582));
    LocalMux I__8473 (
            .O(N__35595),
            .I(N__35579));
    Span4Mux_v I__8472 (
            .O(N__35592),
            .I(N__35576));
    LocalMux I__8471 (
            .O(N__35589),
            .I(N__35573));
    InMux I__8470 (
            .O(N__35588),
            .I(N__35570));
    Span4Mux_v I__8469 (
            .O(N__35585),
            .I(N__35564));
    LocalMux I__8468 (
            .O(N__35582),
            .I(N__35564));
    Span4Mux_h I__8467 (
            .O(N__35579),
            .I(N__35560));
    Span4Mux_v I__8466 (
            .O(N__35576),
            .I(N__35553));
    Span4Mux_v I__8465 (
            .O(N__35573),
            .I(N__35553));
    LocalMux I__8464 (
            .O(N__35570),
            .I(N__35553));
    InMux I__8463 (
            .O(N__35569),
            .I(N__35550));
    Span4Mux_v I__8462 (
            .O(N__35564),
            .I(N__35547));
    InMux I__8461 (
            .O(N__35563),
            .I(N__35544));
    Span4Mux_v I__8460 (
            .O(N__35560),
            .I(N__35539));
    Span4Mux_h I__8459 (
            .O(N__35553),
            .I(N__35539));
    LocalMux I__8458 (
            .O(N__35550),
            .I(N__35536));
    Sp12to4 I__8457 (
            .O(N__35547),
            .I(N__35531));
    LocalMux I__8456 (
            .O(N__35544),
            .I(N__35531));
    Span4Mux_v I__8455 (
            .O(N__35539),
            .I(N__35528));
    Span12Mux_h I__8454 (
            .O(N__35536),
            .I(N__35525));
    Span12Mux_h I__8453 (
            .O(N__35531),
            .I(N__35522));
    Span4Mux_v I__8452 (
            .O(N__35528),
            .I(N__35519));
    Odrv12 I__8451 (
            .O(N__35525),
            .I(port_data_c_0));
    Odrv12 I__8450 (
            .O(N__35522),
            .I(port_data_c_0));
    Odrv4 I__8449 (
            .O(N__35519),
            .I(port_data_c_0));
    InMux I__8448 (
            .O(N__35512),
            .I(N__35508));
    InMux I__8447 (
            .O(N__35511),
            .I(N__35505));
    LocalMux I__8446 (
            .O(N__35508),
            .I(N__35499));
    LocalMux I__8445 (
            .O(N__35505),
            .I(N__35499));
    InMux I__8444 (
            .O(N__35504),
            .I(N__35495));
    Span4Mux_h I__8443 (
            .O(N__35499),
            .I(N__35492));
    InMux I__8442 (
            .O(N__35498),
            .I(N__35488));
    LocalMux I__8441 (
            .O(N__35495),
            .I(N__35485));
    Span4Mux_v I__8440 (
            .O(N__35492),
            .I(N__35482));
    InMux I__8439 (
            .O(N__35491),
            .I(N__35479));
    LocalMux I__8438 (
            .O(N__35488),
            .I(N__35476));
    Span4Mux_v I__8437 (
            .O(N__35485),
            .I(N__35472));
    Span4Mux_v I__8436 (
            .O(N__35482),
            .I(N__35464));
    LocalMux I__8435 (
            .O(N__35479),
            .I(N__35464));
    Span4Mux_v I__8434 (
            .O(N__35476),
            .I(N__35461));
    InMux I__8433 (
            .O(N__35475),
            .I(N__35458));
    Span4Mux_v I__8432 (
            .O(N__35472),
            .I(N__35455));
    InMux I__8431 (
            .O(N__35471),
            .I(N__35450));
    InMux I__8430 (
            .O(N__35470),
            .I(N__35450));
    InMux I__8429 (
            .O(N__35469),
            .I(N__35447));
    Span4Mux_v I__8428 (
            .O(N__35464),
            .I(N__35444));
    Sp12to4 I__8427 (
            .O(N__35461),
            .I(N__35439));
    LocalMux I__8426 (
            .O(N__35458),
            .I(N__35439));
    Sp12to4 I__8425 (
            .O(N__35455),
            .I(N__35432));
    LocalMux I__8424 (
            .O(N__35450),
            .I(N__35432));
    LocalMux I__8423 (
            .O(N__35447),
            .I(N__35432));
    Span4Mux_v I__8422 (
            .O(N__35444),
            .I(N__35429));
    Span12Mux_h I__8421 (
            .O(N__35439),
            .I(N__35426));
    Span12Mux_h I__8420 (
            .O(N__35432),
            .I(N__35423));
    IoSpan4Mux I__8419 (
            .O(N__35429),
            .I(N__35420));
    Odrv12 I__8418 (
            .O(N__35426),
            .I(port_data_c_1));
    Odrv12 I__8417 (
            .O(N__35423),
            .I(port_data_c_1));
    Odrv4 I__8416 (
            .O(N__35420),
            .I(port_data_c_1));
    InMux I__8415 (
            .O(N__35413),
            .I(N__35410));
    LocalMux I__8414 (
            .O(N__35410),
            .I(N__35407));
    Span4Mux_h I__8413 (
            .O(N__35407),
            .I(N__35404));
    Odrv4 I__8412 (
            .O(N__35404),
            .I(\this_ppu.oam_cache.mem_16 ));
    InMux I__8411 (
            .O(N__35401),
            .I(N__35397));
    InMux I__8410 (
            .O(N__35400),
            .I(N__35394));
    LocalMux I__8409 (
            .O(N__35397),
            .I(N__35391));
    LocalMux I__8408 (
            .O(N__35394),
            .I(N__35388));
    Span4Mux_h I__8407 (
            .O(N__35391),
            .I(N__35385));
    Odrv12 I__8406 (
            .O(N__35388),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    Odrv4 I__8405 (
            .O(N__35385),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    InMux I__8404 (
            .O(N__35380),
            .I(N__35377));
    LocalMux I__8403 (
            .O(N__35377),
            .I(N__35374));
    Span4Mux_v I__8402 (
            .O(N__35374),
            .I(N__35371));
    Span4Mux_h I__8401 (
            .O(N__35371),
            .I(N__35368));
    Odrv4 I__8400 (
            .O(N__35368),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__8399 (
            .O(N__35365),
            .I(N__35362));
    LocalMux I__8398 (
            .O(N__35362),
            .I(N__35359));
    Span4Mux_h I__8397 (
            .O(N__35359),
            .I(N__35356));
    Span4Mux_v I__8396 (
            .O(N__35356),
            .I(N__35353));
    Odrv4 I__8395 (
            .O(N__35353),
            .I(M_this_oam_ram_write_data_20));
    InMux I__8394 (
            .O(N__35350),
            .I(N__35347));
    LocalMux I__8393 (
            .O(N__35347),
            .I(N__35344));
    Span4Mux_v I__8392 (
            .O(N__35344),
            .I(N__35341));
    Odrv4 I__8391 (
            .O(N__35341),
            .I(\this_ppu.oam_cache.mem_12 ));
    CascadeMux I__8390 (
            .O(N__35338),
            .I(N__35335));
    InMux I__8389 (
            .O(N__35335),
            .I(N__35329));
    InMux I__8388 (
            .O(N__35334),
            .I(N__35326));
    InMux I__8387 (
            .O(N__35333),
            .I(N__35321));
    InMux I__8386 (
            .O(N__35332),
            .I(N__35318));
    LocalMux I__8385 (
            .O(N__35329),
            .I(N__35315));
    LocalMux I__8384 (
            .O(N__35326),
            .I(N__35312));
    InMux I__8383 (
            .O(N__35325),
            .I(N__35309));
    InMux I__8382 (
            .O(N__35324),
            .I(N__35306));
    LocalMux I__8381 (
            .O(N__35321),
            .I(N__35303));
    LocalMux I__8380 (
            .O(N__35318),
            .I(N__35300));
    Span4Mux_v I__8379 (
            .O(N__35315),
            .I(N__35297));
    Span4Mux_h I__8378 (
            .O(N__35312),
            .I(N__35292));
    LocalMux I__8377 (
            .O(N__35309),
            .I(N__35292));
    LocalMux I__8376 (
            .O(N__35306),
            .I(N__35287));
    Span4Mux_v I__8375 (
            .O(N__35303),
            .I(N__35287));
    Span4Mux_h I__8374 (
            .O(N__35300),
            .I(N__35284));
    Odrv4 I__8373 (
            .O(N__35297),
            .I(\this_ppu.M_hoffset_qZ0Z_2 ));
    Odrv4 I__8372 (
            .O(N__35292),
            .I(\this_ppu.M_hoffset_qZ0Z_2 ));
    Odrv4 I__8371 (
            .O(N__35287),
            .I(\this_ppu.M_hoffset_qZ0Z_2 ));
    Odrv4 I__8370 (
            .O(N__35284),
            .I(\this_ppu.M_hoffset_qZ0Z_2 ));
    CascadeMux I__8369 (
            .O(N__35275),
            .I(N__35272));
    InMux I__8368 (
            .O(N__35272),
            .I(N__35269));
    LocalMux I__8367 (
            .O(N__35269),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0 ));
    InMux I__8366 (
            .O(N__35266),
            .I(N__35263));
    LocalMux I__8365 (
            .O(N__35263),
            .I(N__35260));
    Span4Mux_h I__8364 (
            .O(N__35260),
            .I(N__35257));
    Odrv4 I__8363 (
            .O(N__35257),
            .I(\this_ppu.oam_cache.mem_9 ));
    InMux I__8362 (
            .O(N__35254),
            .I(N__35251));
    LocalMux I__8361 (
            .O(N__35251),
            .I(N__35248));
    Span4Mux_h I__8360 (
            .O(N__35248),
            .I(N__35245));
    Odrv4 I__8359 (
            .O(N__35245),
            .I(\this_ppu.oam_cache.mem_8 ));
    InMux I__8358 (
            .O(N__35242),
            .I(N__35239));
    LocalMux I__8357 (
            .O(N__35239),
            .I(N__35236));
    Span4Mux_h I__8356 (
            .O(N__35236),
            .I(N__35233));
    Odrv4 I__8355 (
            .O(N__35233),
            .I(\this_ppu.oam_cache.mem_13 ));
    InMux I__8354 (
            .O(N__35230),
            .I(N__35221));
    InMux I__8353 (
            .O(N__35229),
            .I(N__35221));
    InMux I__8352 (
            .O(N__35228),
            .I(N__35216));
    InMux I__8351 (
            .O(N__35227),
            .I(N__35216));
    InMux I__8350 (
            .O(N__35226),
            .I(N__35213));
    LocalMux I__8349 (
            .O(N__35221),
            .I(\this_ppu.un1_M_oam_cache_read_data_c4 ));
    LocalMux I__8348 (
            .O(N__35216),
            .I(\this_ppu.un1_M_oam_cache_read_data_c4 ));
    LocalMux I__8347 (
            .O(N__35213),
            .I(\this_ppu.un1_M_oam_cache_read_data_c4 ));
    CascadeMux I__8346 (
            .O(N__35206),
            .I(N__35203));
    CascadeBuf I__8345 (
            .O(N__35203),
            .I(N__35200));
    CascadeMux I__8344 (
            .O(N__35200),
            .I(N__35196));
    CascadeMux I__8343 (
            .O(N__35199),
            .I(N__35193));
    InMux I__8342 (
            .O(N__35196),
            .I(N__35189));
    InMux I__8341 (
            .O(N__35193),
            .I(N__35186));
    InMux I__8340 (
            .O(N__35192),
            .I(N__35183));
    LocalMux I__8339 (
            .O(N__35189),
            .I(N__35179));
    LocalMux I__8338 (
            .O(N__35186),
            .I(N__35175));
    LocalMux I__8337 (
            .O(N__35183),
            .I(N__35171));
    InMux I__8336 (
            .O(N__35182),
            .I(N__35168));
    Span4Mux_h I__8335 (
            .O(N__35179),
            .I(N__35165));
    InMux I__8334 (
            .O(N__35178),
            .I(N__35162));
    Span4Mux_h I__8333 (
            .O(N__35175),
            .I(N__35159));
    InMux I__8332 (
            .O(N__35174),
            .I(N__35156));
    Span4Mux_v I__8331 (
            .O(N__35171),
            .I(N__35151));
    LocalMux I__8330 (
            .O(N__35168),
            .I(N__35151));
    Span4Mux_h I__8329 (
            .O(N__35165),
            .I(N__35148));
    LocalMux I__8328 (
            .O(N__35162),
            .I(N__35141));
    Span4Mux_h I__8327 (
            .O(N__35159),
            .I(N__35141));
    LocalMux I__8326 (
            .O(N__35156),
            .I(N__35141));
    Span4Mux_h I__8325 (
            .O(N__35151),
            .I(N__35136));
    Span4Mux_h I__8324 (
            .O(N__35148),
            .I(N__35136));
    Span4Mux_v I__8323 (
            .O(N__35141),
            .I(N__35133));
    Span4Mux_v I__8322 (
            .O(N__35136),
            .I(N__35130));
    Odrv4 I__8321 (
            .O(N__35133),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__8320 (
            .O(N__35130),
            .I(M_this_ppu_map_addr_2));
    InMux I__8319 (
            .O(N__35125),
            .I(N__35121));
    InMux I__8318 (
            .O(N__35124),
            .I(N__35118));
    LocalMux I__8317 (
            .O(N__35121),
            .I(N__35112));
    LocalMux I__8316 (
            .O(N__35118),
            .I(N__35112));
    InMux I__8315 (
            .O(N__35117),
            .I(N__35109));
    Span4Mux_h I__8314 (
            .O(N__35112),
            .I(N__35103));
    LocalMux I__8313 (
            .O(N__35109),
            .I(N__35100));
    InMux I__8312 (
            .O(N__35108),
            .I(N__35097));
    InMux I__8311 (
            .O(N__35107),
            .I(N__35094));
    InMux I__8310 (
            .O(N__35106),
            .I(N__35091));
    Odrv4 I__8309 (
            .O(N__35103),
            .I(\this_ppu.un1_M_hoffset_q_8 ));
    Odrv4 I__8308 (
            .O(N__35100),
            .I(\this_ppu.un1_M_hoffset_q_8 ));
    LocalMux I__8307 (
            .O(N__35097),
            .I(\this_ppu.un1_M_hoffset_q_8 ));
    LocalMux I__8306 (
            .O(N__35094),
            .I(\this_ppu.un1_M_hoffset_q_8 ));
    LocalMux I__8305 (
            .O(N__35091),
            .I(\this_ppu.un1_M_hoffset_q_8 ));
    CascadeMux I__8304 (
            .O(N__35080),
            .I(\this_ppu.un1_M_oam_cache_read_data_c4_cascade_ ));
    InMux I__8303 (
            .O(N__35077),
            .I(N__35074));
    LocalMux I__8302 (
            .O(N__35074),
            .I(N__35069));
    CascadeMux I__8301 (
            .O(N__35073),
            .I(N__35066));
    InMux I__8300 (
            .O(N__35072),
            .I(N__35058));
    Span4Mux_h I__8299 (
            .O(N__35069),
            .I(N__35055));
    InMux I__8298 (
            .O(N__35066),
            .I(N__35050));
    InMux I__8297 (
            .O(N__35065),
            .I(N__35050));
    InMux I__8296 (
            .O(N__35064),
            .I(N__35047));
    InMux I__8295 (
            .O(N__35063),
            .I(N__35042));
    InMux I__8294 (
            .O(N__35062),
            .I(N__35042));
    InMux I__8293 (
            .O(N__35061),
            .I(N__35039));
    LocalMux I__8292 (
            .O(N__35058),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    Odrv4 I__8291 (
            .O(N__35055),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    LocalMux I__8290 (
            .O(N__35050),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    LocalMux I__8289 (
            .O(N__35047),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    LocalMux I__8288 (
            .O(N__35042),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    LocalMux I__8287 (
            .O(N__35039),
            .I(\this_ppu.un1_M_hoffset_q_7 ));
    InMux I__8286 (
            .O(N__35026),
            .I(N__35023));
    LocalMux I__8285 (
            .O(N__35023),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0 ));
    InMux I__8284 (
            .O(N__35020),
            .I(N__35017));
    LocalMux I__8283 (
            .O(N__35017),
            .I(N__35014));
    Span4Mux_h I__8282 (
            .O(N__35014),
            .I(N__35010));
    InMux I__8281 (
            .O(N__35013),
            .I(N__35007));
    Odrv4 I__8280 (
            .O(N__35010),
            .I(\this_ppu.read_data_RNI80ET_11 ));
    LocalMux I__8279 (
            .O(N__35007),
            .I(\this_ppu.read_data_RNI80ET_11 ));
    InMux I__8278 (
            .O(N__35002),
            .I(N__34999));
    LocalMux I__8277 (
            .O(N__34999),
            .I(N__34996));
    Span4Mux_h I__8276 (
            .O(N__34996),
            .I(N__34993));
    Odrv4 I__8275 (
            .O(N__34993),
            .I(M_this_oam_ram_read_data_11));
    InMux I__8274 (
            .O(N__34990),
            .I(N__34987));
    LocalMux I__8273 (
            .O(N__34987),
            .I(N__34984));
    Odrv4 I__8272 (
            .O(N__34984),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_11 ));
    InMux I__8271 (
            .O(N__34981),
            .I(N__34978));
    LocalMux I__8270 (
            .O(N__34978),
            .I(N__34972));
    InMux I__8269 (
            .O(N__34977),
            .I(N__34969));
    InMux I__8268 (
            .O(N__34976),
            .I(N__34963));
    InMux I__8267 (
            .O(N__34975),
            .I(N__34959));
    Span4Mux_v I__8266 (
            .O(N__34972),
            .I(N__34951));
    LocalMux I__8265 (
            .O(N__34969),
            .I(N__34951));
    InMux I__8264 (
            .O(N__34968),
            .I(N__34948));
    InMux I__8263 (
            .O(N__34967),
            .I(N__34945));
    InMux I__8262 (
            .O(N__34966),
            .I(N__34942));
    LocalMux I__8261 (
            .O(N__34963),
            .I(N__34937));
    InMux I__8260 (
            .O(N__34962),
            .I(N__34934));
    LocalMux I__8259 (
            .O(N__34959),
            .I(N__34931));
    InMux I__8258 (
            .O(N__34958),
            .I(N__34924));
    InMux I__8257 (
            .O(N__34957),
            .I(N__34924));
    InMux I__8256 (
            .O(N__34956),
            .I(N__34924));
    Span4Mux_v I__8255 (
            .O(N__34951),
            .I(N__34918));
    LocalMux I__8254 (
            .O(N__34948),
            .I(N__34918));
    LocalMux I__8253 (
            .O(N__34945),
            .I(N__34913));
    LocalMux I__8252 (
            .O(N__34942),
            .I(N__34913));
    InMux I__8251 (
            .O(N__34941),
            .I(N__34908));
    InMux I__8250 (
            .O(N__34940),
            .I(N__34908));
    Span4Mux_v I__8249 (
            .O(N__34937),
            .I(N__34903));
    LocalMux I__8248 (
            .O(N__34934),
            .I(N__34903));
    Span4Mux_v I__8247 (
            .O(N__34931),
            .I(N__34898));
    LocalMux I__8246 (
            .O(N__34924),
            .I(N__34898));
    InMux I__8245 (
            .O(N__34923),
            .I(N__34895));
    Span4Mux_v I__8244 (
            .O(N__34918),
            .I(N__34892));
    Span4Mux_h I__8243 (
            .O(N__34913),
            .I(N__34889));
    LocalMux I__8242 (
            .O(N__34908),
            .I(N__34886));
    Span4Mux_v I__8241 (
            .O(N__34903),
            .I(N__34883));
    Span4Mux_h I__8240 (
            .O(N__34898),
            .I(N__34880));
    LocalMux I__8239 (
            .O(N__34895),
            .I(N__34877));
    Span4Mux_h I__8238 (
            .O(N__34892),
            .I(N__34874));
    Span4Mux_v I__8237 (
            .O(N__34889),
            .I(N__34869));
    Span4Mux_v I__8236 (
            .O(N__34886),
            .I(N__34869));
    Odrv4 I__8235 (
            .O(N__34883),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv4 I__8234 (
            .O(N__34880),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv12 I__8233 (
            .O(N__34877),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv4 I__8232 (
            .O(N__34874),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv4 I__8231 (
            .O(N__34869),
            .I(\this_ppu.M_state_q_inv_1 ));
    InMux I__8230 (
            .O(N__34858),
            .I(N__34854));
    CascadeMux I__8229 (
            .O(N__34857),
            .I(N__34851));
    LocalMux I__8228 (
            .O(N__34854),
            .I(N__34847));
    InMux I__8227 (
            .O(N__34851),
            .I(N__34844));
    InMux I__8226 (
            .O(N__34850),
            .I(N__34840));
    Span4Mux_h I__8225 (
            .O(N__34847),
            .I(N__34834));
    LocalMux I__8224 (
            .O(N__34844),
            .I(N__34834));
    InMux I__8223 (
            .O(N__34843),
            .I(N__34831));
    LocalMux I__8222 (
            .O(N__34840),
            .I(N__34828));
    InMux I__8221 (
            .O(N__34839),
            .I(N__34825));
    Span4Mux_v I__8220 (
            .O(N__34834),
            .I(N__34822));
    LocalMux I__8219 (
            .O(N__34831),
            .I(N__34817));
    Span4Mux_v I__8218 (
            .O(N__34828),
            .I(N__34817));
    LocalMux I__8217 (
            .O(N__34825),
            .I(\this_ppu.vspr ));
    Odrv4 I__8216 (
            .O(N__34822),
            .I(\this_ppu.vspr ));
    Odrv4 I__8215 (
            .O(N__34817),
            .I(\this_ppu.vspr ));
    CascadeMux I__8214 (
            .O(N__34810),
            .I(N__34804));
    CascadeMux I__8213 (
            .O(N__34809),
            .I(N__34801));
    CascadeMux I__8212 (
            .O(N__34808),
            .I(N__34789));
    CascadeMux I__8211 (
            .O(N__34807),
            .I(N__34786));
    InMux I__8210 (
            .O(N__34804),
            .I(N__34782));
    InMux I__8209 (
            .O(N__34801),
            .I(N__34779));
    CascadeMux I__8208 (
            .O(N__34800),
            .I(N__34776));
    CascadeMux I__8207 (
            .O(N__34799),
            .I(N__34773));
    CascadeMux I__8206 (
            .O(N__34798),
            .I(N__34770));
    CascadeMux I__8205 (
            .O(N__34797),
            .I(N__34767));
    CascadeMux I__8204 (
            .O(N__34796),
            .I(N__34764));
    CascadeMux I__8203 (
            .O(N__34795),
            .I(N__34761));
    CascadeMux I__8202 (
            .O(N__34794),
            .I(N__34757));
    CascadeMux I__8201 (
            .O(N__34793),
            .I(N__34754));
    CascadeMux I__8200 (
            .O(N__34792),
            .I(N__34751));
    InMux I__8199 (
            .O(N__34789),
            .I(N__34748));
    InMux I__8198 (
            .O(N__34786),
            .I(N__34745));
    CascadeMux I__8197 (
            .O(N__34785),
            .I(N__34742));
    LocalMux I__8196 (
            .O(N__34782),
            .I(N__34737));
    LocalMux I__8195 (
            .O(N__34779),
            .I(N__34737));
    InMux I__8194 (
            .O(N__34776),
            .I(N__34734));
    InMux I__8193 (
            .O(N__34773),
            .I(N__34731));
    InMux I__8192 (
            .O(N__34770),
            .I(N__34728));
    InMux I__8191 (
            .O(N__34767),
            .I(N__34724));
    InMux I__8190 (
            .O(N__34764),
            .I(N__34721));
    InMux I__8189 (
            .O(N__34761),
            .I(N__34718));
    CascadeMux I__8188 (
            .O(N__34760),
            .I(N__34715));
    InMux I__8187 (
            .O(N__34757),
            .I(N__34712));
    InMux I__8186 (
            .O(N__34754),
            .I(N__34709));
    InMux I__8185 (
            .O(N__34751),
            .I(N__34706));
    LocalMux I__8184 (
            .O(N__34748),
            .I(N__34703));
    LocalMux I__8183 (
            .O(N__34745),
            .I(N__34700));
    InMux I__8182 (
            .O(N__34742),
            .I(N__34697));
    Span4Mux_v I__8181 (
            .O(N__34737),
            .I(N__34690));
    LocalMux I__8180 (
            .O(N__34734),
            .I(N__34690));
    LocalMux I__8179 (
            .O(N__34731),
            .I(N__34690));
    LocalMux I__8178 (
            .O(N__34728),
            .I(N__34687));
    CascadeMux I__8177 (
            .O(N__34727),
            .I(N__34684));
    LocalMux I__8176 (
            .O(N__34724),
            .I(N__34679));
    LocalMux I__8175 (
            .O(N__34721),
            .I(N__34679));
    LocalMux I__8174 (
            .O(N__34718),
            .I(N__34676));
    InMux I__8173 (
            .O(N__34715),
            .I(N__34673));
    LocalMux I__8172 (
            .O(N__34712),
            .I(N__34670));
    LocalMux I__8171 (
            .O(N__34709),
            .I(N__34665));
    LocalMux I__8170 (
            .O(N__34706),
            .I(N__34665));
    Span4Mux_v I__8169 (
            .O(N__34703),
            .I(N__34660));
    Span4Mux_s1_v I__8168 (
            .O(N__34700),
            .I(N__34660));
    LocalMux I__8167 (
            .O(N__34697),
            .I(N__34657));
    Span4Mux_v I__8166 (
            .O(N__34690),
            .I(N__34652));
    Span4Mux_v I__8165 (
            .O(N__34687),
            .I(N__34652));
    InMux I__8164 (
            .O(N__34684),
            .I(N__34649));
    Span4Mux_v I__8163 (
            .O(N__34679),
            .I(N__34644));
    Span4Mux_v I__8162 (
            .O(N__34676),
            .I(N__34644));
    LocalMux I__8161 (
            .O(N__34673),
            .I(N__34641));
    Span4Mux_v I__8160 (
            .O(N__34670),
            .I(N__34634));
    Span4Mux_v I__8159 (
            .O(N__34665),
            .I(N__34634));
    Span4Mux_v I__8158 (
            .O(N__34660),
            .I(N__34634));
    Span4Mux_v I__8157 (
            .O(N__34657),
            .I(N__34631));
    Sp12to4 I__8156 (
            .O(N__34652),
            .I(N__34628));
    LocalMux I__8155 (
            .O(N__34649),
            .I(N__34625));
    Span4Mux_h I__8154 (
            .O(N__34644),
            .I(N__34622));
    Span4Mux_v I__8153 (
            .O(N__34641),
            .I(N__34619));
    Sp12to4 I__8152 (
            .O(N__34634),
            .I(N__34616));
    Sp12to4 I__8151 (
            .O(N__34631),
            .I(N__34613));
    Span12Mux_h I__8150 (
            .O(N__34628),
            .I(N__34610));
    Span4Mux_v I__8149 (
            .O(N__34625),
            .I(N__34603));
    Span4Mux_v I__8148 (
            .O(N__34622),
            .I(N__34603));
    Span4Mux_v I__8147 (
            .O(N__34619),
            .I(N__34603));
    Span12Mux_s9_h I__8146 (
            .O(N__34616),
            .I(N__34600));
    Span12Mux_h I__8145 (
            .O(N__34613),
            .I(N__34595));
    Span12Mux_v I__8144 (
            .O(N__34610),
            .I(N__34595));
    Odrv4 I__8143 (
            .O(N__34603),
            .I(M_this_ppu_spr_addr_3));
    Odrv12 I__8142 (
            .O(N__34600),
            .I(M_this_ppu_spr_addr_3));
    Odrv12 I__8141 (
            .O(N__34595),
            .I(M_this_ppu_spr_addr_3));
    InMux I__8140 (
            .O(N__34588),
            .I(N__34585));
    LocalMux I__8139 (
            .O(N__34585),
            .I(N__34582));
    Span4Mux_h I__8138 (
            .O(N__34582),
            .I(N__34579));
    Odrv4 I__8137 (
            .O(N__34579),
            .I(\this_ppu.oam_cache.mem_15 ));
    InMux I__8136 (
            .O(N__34576),
            .I(N__34573));
    LocalMux I__8135 (
            .O(N__34573),
            .I(N__34570));
    Span4Mux_h I__8134 (
            .O(N__34570),
            .I(N__34567));
    Odrv4 I__8133 (
            .O(N__34567),
            .I(\this_ppu.oam_cache.mem_14 ));
    InMux I__8132 (
            .O(N__34564),
            .I(N__34561));
    LocalMux I__8131 (
            .O(N__34561),
            .I(N__34555));
    InMux I__8130 (
            .O(N__34560),
            .I(N__34547));
    InMux I__8129 (
            .O(N__34559),
            .I(N__34547));
    InMux I__8128 (
            .O(N__34558),
            .I(N__34547));
    Span4Mux_v I__8127 (
            .O(N__34555),
            .I(N__34544));
    InMux I__8126 (
            .O(N__34554),
            .I(N__34541));
    LocalMux I__8125 (
            .O(N__34547),
            .I(N__34538));
    Span4Mux_v I__8124 (
            .O(N__34544),
            .I(N__34535));
    LocalMux I__8123 (
            .O(N__34541),
            .I(N__34532));
    Span4Mux_h I__8122 (
            .O(N__34538),
            .I(N__34529));
    Span4Mux_v I__8121 (
            .O(N__34535),
            .I(N__34526));
    Span4Mux_h I__8120 (
            .O(N__34532),
            .I(N__34521));
    Span4Mux_v I__8119 (
            .O(N__34529),
            .I(N__34521));
    Odrv4 I__8118 (
            .O(N__34526),
            .I(M_this_oam_ram_read_data_22));
    Odrv4 I__8117 (
            .O(N__34521),
            .I(M_this_oam_ram_read_data_22));
    InMux I__8116 (
            .O(N__34516),
            .I(N__34513));
    LocalMux I__8115 (
            .O(N__34513),
            .I(N__34510));
    Span4Mux_v I__8114 (
            .O(N__34510),
            .I(N__34507));
    Span4Mux_v I__8113 (
            .O(N__34507),
            .I(N__34504));
    Odrv4 I__8112 (
            .O(N__34504),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_22 ));
    InMux I__8111 (
            .O(N__34501),
            .I(N__34496));
    CascadeMux I__8110 (
            .O(N__34500),
            .I(N__34492));
    CascadeMux I__8109 (
            .O(N__34499),
            .I(N__34489));
    LocalMux I__8108 (
            .O(N__34496),
            .I(N__34485));
    InMux I__8107 (
            .O(N__34495),
            .I(N__34475));
    InMux I__8106 (
            .O(N__34492),
            .I(N__34475));
    InMux I__8105 (
            .O(N__34489),
            .I(N__34475));
    InMux I__8104 (
            .O(N__34488),
            .I(N__34475));
    Span4Mux_h I__8103 (
            .O(N__34485),
            .I(N__34472));
    InMux I__8102 (
            .O(N__34484),
            .I(N__34469));
    LocalMux I__8101 (
            .O(N__34475),
            .I(N__34466));
    Span4Mux_v I__8100 (
            .O(N__34472),
            .I(N__34463));
    LocalMux I__8099 (
            .O(N__34469),
            .I(N__34460));
    Span4Mux_h I__8098 (
            .O(N__34466),
            .I(N__34457));
    Span4Mux_v I__8097 (
            .O(N__34463),
            .I(N__34454));
    Span4Mux_h I__8096 (
            .O(N__34460),
            .I(N__34449));
    Span4Mux_v I__8095 (
            .O(N__34457),
            .I(N__34449));
    Odrv4 I__8094 (
            .O(N__34454),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__8093 (
            .O(N__34449),
            .I(M_this_oam_ram_read_data_21));
    InMux I__8092 (
            .O(N__34444),
            .I(N__34441));
    LocalMux I__8091 (
            .O(N__34441),
            .I(N__34438));
    Span4Mux_h I__8090 (
            .O(N__34438),
            .I(N__34435));
    Span4Mux_v I__8089 (
            .O(N__34435),
            .I(N__34432));
    Odrv4 I__8088 (
            .O(N__34432),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_21 ));
    CascadeMux I__8087 (
            .O(N__34429),
            .I(N__34424));
    InMux I__8086 (
            .O(N__34428),
            .I(N__34420));
    InMux I__8085 (
            .O(N__34427),
            .I(N__34417));
    InMux I__8084 (
            .O(N__34424),
            .I(N__34414));
    CascadeMux I__8083 (
            .O(N__34423),
            .I(N__34411));
    LocalMux I__8082 (
            .O(N__34420),
            .I(N__34406));
    LocalMux I__8081 (
            .O(N__34417),
            .I(N__34406));
    LocalMux I__8080 (
            .O(N__34414),
            .I(N__34403));
    InMux I__8079 (
            .O(N__34411),
            .I(N__34400));
    Odrv4 I__8078 (
            .O(N__34406),
            .I(\this_ppu.un1_M_hoffset_q_9 ));
    Odrv4 I__8077 (
            .O(N__34403),
            .I(\this_ppu.un1_M_hoffset_q_9 ));
    LocalMux I__8076 (
            .O(N__34400),
            .I(\this_ppu.un1_M_hoffset_q_9 ));
    InMux I__8075 (
            .O(N__34393),
            .I(N__34387));
    InMux I__8074 (
            .O(N__34392),
            .I(N__34387));
    LocalMux I__8073 (
            .O(N__34387),
            .I(N__34381));
    InMux I__8072 (
            .O(N__34386),
            .I(N__34374));
    InMux I__8071 (
            .O(N__34385),
            .I(N__34374));
    InMux I__8070 (
            .O(N__34384),
            .I(N__34374));
    Odrv4 I__8069 (
            .O(N__34381),
            .I(\this_ppu.un1_M_oam_cache_read_data_c7 ));
    LocalMux I__8068 (
            .O(N__34374),
            .I(\this_ppu.un1_M_oam_cache_read_data_c7 ));
    CascadeMux I__8067 (
            .O(N__34369),
            .I(N__34363));
    CascadeMux I__8066 (
            .O(N__34368),
            .I(N__34360));
    InMux I__8065 (
            .O(N__34367),
            .I(N__34355));
    InMux I__8064 (
            .O(N__34366),
            .I(N__34355));
    InMux I__8063 (
            .O(N__34363),
            .I(N__34351));
    InMux I__8062 (
            .O(N__34360),
            .I(N__34348));
    LocalMux I__8061 (
            .O(N__34355),
            .I(N__34345));
    InMux I__8060 (
            .O(N__34354),
            .I(N__34339));
    LocalMux I__8059 (
            .O(N__34351),
            .I(N__34336));
    LocalMux I__8058 (
            .O(N__34348),
            .I(N__34333));
    Span4Mux_h I__8057 (
            .O(N__34345),
            .I(N__34330));
    InMux I__8056 (
            .O(N__34344),
            .I(N__34325));
    InMux I__8055 (
            .O(N__34343),
            .I(N__34325));
    InMux I__8054 (
            .O(N__34342),
            .I(N__34322));
    LocalMux I__8053 (
            .O(N__34339),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    Odrv4 I__8052 (
            .O(N__34336),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    Odrv12 I__8051 (
            .O(N__34333),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    Odrv4 I__8050 (
            .O(N__34330),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    LocalMux I__8049 (
            .O(N__34325),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    LocalMux I__8048 (
            .O(N__34322),
            .I(\this_ppu.un1_M_hoffset_q_10 ));
    CascadeMux I__8047 (
            .O(N__34309),
            .I(\this_ppu.un1_M_oam_cache_read_data_c7_cascade_ ));
    CascadeMux I__8046 (
            .O(N__34306),
            .I(N__34303));
    CascadeBuf I__8045 (
            .O(N__34303),
            .I(N__34297));
    CascadeMux I__8044 (
            .O(N__34302),
            .I(N__34293));
    InMux I__8043 (
            .O(N__34301),
            .I(N__34290));
    InMux I__8042 (
            .O(N__34300),
            .I(N__34287));
    CascadeMux I__8041 (
            .O(N__34297),
            .I(N__34283));
    InMux I__8040 (
            .O(N__34296),
            .I(N__34280));
    InMux I__8039 (
            .O(N__34293),
            .I(N__34277));
    LocalMux I__8038 (
            .O(N__34290),
            .I(N__34272));
    LocalMux I__8037 (
            .O(N__34287),
            .I(N__34272));
    InMux I__8036 (
            .O(N__34286),
            .I(N__34269));
    InMux I__8035 (
            .O(N__34283),
            .I(N__34266));
    LocalMux I__8034 (
            .O(N__34280),
            .I(N__34261));
    LocalMux I__8033 (
            .O(N__34277),
            .I(N__34261));
    Span4Mux_v I__8032 (
            .O(N__34272),
            .I(N__34256));
    LocalMux I__8031 (
            .O(N__34269),
            .I(N__34256));
    LocalMux I__8030 (
            .O(N__34266),
            .I(N__34253));
    Span4Mux_h I__8029 (
            .O(N__34261),
            .I(N__34250));
    Span4Mux_h I__8028 (
            .O(N__34256),
            .I(N__34247));
    Span12Mux_v I__8027 (
            .O(N__34253),
            .I(N__34244));
    Odrv4 I__8026 (
            .O(N__34250),
            .I(M_this_ppu_map_addr_4));
    Odrv4 I__8025 (
            .O(N__34247),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__8024 (
            .O(N__34244),
            .I(M_this_ppu_map_addr_4));
    CascadeMux I__8023 (
            .O(N__34237),
            .I(N__34234));
    InMux I__8022 (
            .O(N__34234),
            .I(N__34231));
    LocalMux I__8021 (
            .O(N__34231),
            .I(N__34228));
    Odrv4 I__8020 (
            .O(N__34228),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0 ));
    CascadeMux I__8019 (
            .O(N__34225),
            .I(N__34222));
    InMux I__8018 (
            .O(N__34222),
            .I(N__34219));
    LocalMux I__8017 (
            .O(N__34219),
            .I(N__34216));
    Odrv12 I__8016 (
            .O(N__34216),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0 ));
    CEMux I__8015 (
            .O(N__34213),
            .I(N__34209));
    CEMux I__8014 (
            .O(N__34212),
            .I(N__34206));
    LocalMux I__8013 (
            .O(N__34209),
            .I(N__34203));
    LocalMux I__8012 (
            .O(N__34206),
            .I(N__34200));
    Span4Mux_h I__8011 (
            .O(N__34203),
            .I(N__34197));
    Span12Mux_s10_v I__8010 (
            .O(N__34200),
            .I(N__34194));
    Span4Mux_v I__8009 (
            .O(N__34197),
            .I(N__34191));
    Odrv12 I__8008 (
            .O(N__34194),
            .I(\this_spr_ram.mem_WE_0 ));
    Odrv4 I__8007 (
            .O(N__34191),
            .I(\this_spr_ram.mem_WE_0 ));
    InMux I__8006 (
            .O(N__34186),
            .I(N__34183));
    LocalMux I__8005 (
            .O(N__34183),
            .I(N__34180));
    Span4Mux_h I__8004 (
            .O(N__34180),
            .I(N__34177));
    Span4Mux_v I__8003 (
            .O(N__34177),
            .I(N__34174));
    Odrv4 I__8002 (
            .O(N__34174),
            .I(\this_ppu.oam_cache.mem_7 ));
    InMux I__8001 (
            .O(N__34171),
            .I(N__34168));
    LocalMux I__8000 (
            .O(N__34168),
            .I(N__34165));
    Span4Mux_h I__7999 (
            .O(N__34165),
            .I(N__34162));
    Odrv4 I__7998 (
            .O(N__34162),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_7 ));
    CascadeMux I__7997 (
            .O(N__34159),
            .I(N__34155));
    InMux I__7996 (
            .O(N__34158),
            .I(N__34151));
    InMux I__7995 (
            .O(N__34155),
            .I(N__34148));
    CascadeMux I__7994 (
            .O(N__34154),
            .I(N__34145));
    LocalMux I__7993 (
            .O(N__34151),
            .I(N__34139));
    LocalMux I__7992 (
            .O(N__34148),
            .I(N__34139));
    InMux I__7991 (
            .O(N__34145),
            .I(N__34136));
    CascadeMux I__7990 (
            .O(N__34144),
            .I(N__34131));
    Span4Mux_v I__7989 (
            .O(N__34139),
            .I(N__34128));
    LocalMux I__7988 (
            .O(N__34136),
            .I(N__34125));
    InMux I__7987 (
            .O(N__34135),
            .I(N__34121));
    InMux I__7986 (
            .O(N__34134),
            .I(N__34118));
    InMux I__7985 (
            .O(N__34131),
            .I(N__34115));
    Span4Mux_h I__7984 (
            .O(N__34128),
            .I(N__34110));
    Span4Mux_h I__7983 (
            .O(N__34125),
            .I(N__34110));
    InMux I__7982 (
            .O(N__34124),
            .I(N__34107));
    LocalMux I__7981 (
            .O(N__34121),
            .I(\this_ppu.hspr ));
    LocalMux I__7980 (
            .O(N__34118),
            .I(\this_ppu.hspr ));
    LocalMux I__7979 (
            .O(N__34115),
            .I(\this_ppu.hspr ));
    Odrv4 I__7978 (
            .O(N__34110),
            .I(\this_ppu.hspr ));
    LocalMux I__7977 (
            .O(N__34107),
            .I(\this_ppu.hspr ));
    CascadeMux I__7976 (
            .O(N__34096),
            .I(N__34092));
    CascadeMux I__7975 (
            .O(N__34095),
            .I(N__34089));
    InMux I__7974 (
            .O(N__34092),
            .I(N__34082));
    InMux I__7973 (
            .O(N__34089),
            .I(N__34079));
    CascadeMux I__7972 (
            .O(N__34088),
            .I(N__34076));
    CascadeMux I__7971 (
            .O(N__34087),
            .I(N__34073));
    CascadeMux I__7970 (
            .O(N__34086),
            .I(N__34069));
    CascadeMux I__7969 (
            .O(N__34085),
            .I(N__34066));
    LocalMux I__7968 (
            .O(N__34082),
            .I(N__34059));
    LocalMux I__7967 (
            .O(N__34079),
            .I(N__34059));
    InMux I__7966 (
            .O(N__34076),
            .I(N__34056));
    InMux I__7965 (
            .O(N__34073),
            .I(N__34053));
    CascadeMux I__7964 (
            .O(N__34072),
            .I(N__34050));
    InMux I__7963 (
            .O(N__34069),
            .I(N__34047));
    InMux I__7962 (
            .O(N__34066),
            .I(N__34044));
    CascadeMux I__7961 (
            .O(N__34065),
            .I(N__34041));
    CascadeMux I__7960 (
            .O(N__34064),
            .I(N__34038));
    Span4Mux_v I__7959 (
            .O(N__34059),
            .I(N__34030));
    LocalMux I__7958 (
            .O(N__34056),
            .I(N__34030));
    LocalMux I__7957 (
            .O(N__34053),
            .I(N__34030));
    InMux I__7956 (
            .O(N__34050),
            .I(N__34027));
    LocalMux I__7955 (
            .O(N__34047),
            .I(N__34022));
    LocalMux I__7954 (
            .O(N__34044),
            .I(N__34022));
    InMux I__7953 (
            .O(N__34041),
            .I(N__34019));
    InMux I__7952 (
            .O(N__34038),
            .I(N__34016));
    CascadeMux I__7951 (
            .O(N__34037),
            .I(N__34013));
    Span4Mux_v I__7950 (
            .O(N__34030),
            .I(N__34006));
    LocalMux I__7949 (
            .O(N__34027),
            .I(N__34006));
    Span4Mux_s2_v I__7948 (
            .O(N__34022),
            .I(N__34001));
    LocalMux I__7947 (
            .O(N__34019),
            .I(N__34001));
    LocalMux I__7946 (
            .O(N__34016),
            .I(N__33998));
    InMux I__7945 (
            .O(N__34013),
            .I(N__33995));
    CascadeMux I__7944 (
            .O(N__34012),
            .I(N__33990));
    CascadeMux I__7943 (
            .O(N__34011),
            .I(N__33985));
    Span4Mux_v I__7942 (
            .O(N__34006),
            .I(N__33982));
    Span4Mux_v I__7941 (
            .O(N__34001),
            .I(N__33975));
    Span4Mux_h I__7940 (
            .O(N__33998),
            .I(N__33975));
    LocalMux I__7939 (
            .O(N__33995),
            .I(N__33975));
    CascadeMux I__7938 (
            .O(N__33994),
            .I(N__33972));
    CascadeMux I__7937 (
            .O(N__33993),
            .I(N__33969));
    InMux I__7936 (
            .O(N__33990),
            .I(N__33966));
    CascadeMux I__7935 (
            .O(N__33989),
            .I(N__33963));
    CascadeMux I__7934 (
            .O(N__33988),
            .I(N__33960));
    InMux I__7933 (
            .O(N__33985),
            .I(N__33957));
    Span4Mux_h I__7932 (
            .O(N__33982),
            .I(N__33954));
    Span4Mux_v I__7931 (
            .O(N__33975),
            .I(N__33951));
    InMux I__7930 (
            .O(N__33972),
            .I(N__33948));
    InMux I__7929 (
            .O(N__33969),
            .I(N__33945));
    LocalMux I__7928 (
            .O(N__33966),
            .I(N__33942));
    InMux I__7927 (
            .O(N__33963),
            .I(N__33939));
    InMux I__7926 (
            .O(N__33960),
            .I(N__33936));
    LocalMux I__7925 (
            .O(N__33957),
            .I(N__33933));
    Span4Mux_h I__7924 (
            .O(N__33954),
            .I(N__33930));
    Span4Mux_v I__7923 (
            .O(N__33951),
            .I(N__33923));
    LocalMux I__7922 (
            .O(N__33948),
            .I(N__33923));
    LocalMux I__7921 (
            .O(N__33945),
            .I(N__33923));
    Span4Mux_h I__7920 (
            .O(N__33942),
            .I(N__33918));
    LocalMux I__7919 (
            .O(N__33939),
            .I(N__33918));
    LocalMux I__7918 (
            .O(N__33936),
            .I(N__33915));
    Span12Mux_h I__7917 (
            .O(N__33933),
            .I(N__33912));
    Span4Mux_h I__7916 (
            .O(N__33930),
            .I(N__33903));
    Span4Mux_v I__7915 (
            .O(N__33923),
            .I(N__33903));
    Span4Mux_v I__7914 (
            .O(N__33918),
            .I(N__33903));
    Span4Mux_h I__7913 (
            .O(N__33915),
            .I(N__33903));
    Odrv12 I__7912 (
            .O(N__33912),
            .I(M_this_ppu_spr_addr_0));
    Odrv4 I__7911 (
            .O(N__33903),
            .I(M_this_ppu_spr_addr_0));
    InMux I__7910 (
            .O(N__33898),
            .I(N__33895));
    LocalMux I__7909 (
            .O(N__33895),
            .I(N__33891));
    InMux I__7908 (
            .O(N__33894),
            .I(N__33888));
    Span4Mux_h I__7907 (
            .O(N__33891),
            .I(N__33884));
    LocalMux I__7906 (
            .O(N__33888),
            .I(N__33881));
    InMux I__7905 (
            .O(N__33887),
            .I(N__33878));
    Span4Mux_v I__7904 (
            .O(N__33884),
            .I(N__33871));
    Span4Mux_h I__7903 (
            .O(N__33881),
            .I(N__33871));
    LocalMux I__7902 (
            .O(N__33878),
            .I(N__33868));
    InMux I__7901 (
            .O(N__33877),
            .I(N__33865));
    InMux I__7900 (
            .O(N__33876),
            .I(N__33860));
    Span4Mux_h I__7899 (
            .O(N__33871),
            .I(N__33857));
    Span4Mux_h I__7898 (
            .O(N__33868),
            .I(N__33854));
    LocalMux I__7897 (
            .O(N__33865),
            .I(N__33851));
    InMux I__7896 (
            .O(N__33864),
            .I(N__33848));
    InMux I__7895 (
            .O(N__33863),
            .I(N__33845));
    LocalMux I__7894 (
            .O(N__33860),
            .I(N__33841));
    Span4Mux_h I__7893 (
            .O(N__33857),
            .I(N__33838));
    Span4Mux_v I__7892 (
            .O(N__33854),
            .I(N__33833));
    Span4Mux_h I__7891 (
            .O(N__33851),
            .I(N__33833));
    LocalMux I__7890 (
            .O(N__33848),
            .I(N__33830));
    LocalMux I__7889 (
            .O(N__33845),
            .I(N__33827));
    InMux I__7888 (
            .O(N__33844),
            .I(N__33824));
    Span12Mux_h I__7887 (
            .O(N__33841),
            .I(N__33821));
    Span4Mux_h I__7886 (
            .O(N__33838),
            .I(N__33814));
    Span4Mux_v I__7885 (
            .O(N__33833),
            .I(N__33814));
    Span4Mux_h I__7884 (
            .O(N__33830),
            .I(N__33814));
    Span4Mux_v I__7883 (
            .O(N__33827),
            .I(N__33809));
    LocalMux I__7882 (
            .O(N__33824),
            .I(N__33809));
    Odrv12 I__7881 (
            .O(N__33821),
            .I(M_this_spr_ram_write_data_0));
    Odrv4 I__7880 (
            .O(N__33814),
            .I(M_this_spr_ram_write_data_0));
    Odrv4 I__7879 (
            .O(N__33809),
            .I(M_this_spr_ram_write_data_0));
    InMux I__7878 (
            .O(N__33802),
            .I(N__33799));
    LocalMux I__7877 (
            .O(N__33799),
            .I(\this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2 ));
    InMux I__7876 (
            .O(N__33796),
            .I(N__33793));
    LocalMux I__7875 (
            .O(N__33793),
            .I(\this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3 ));
    InMux I__7874 (
            .O(N__33790),
            .I(N__33786));
    InMux I__7873 (
            .O(N__33789),
            .I(N__33783));
    LocalMux I__7872 (
            .O(N__33786),
            .I(N__33780));
    LocalMux I__7871 (
            .O(N__33783),
            .I(N__33775));
    Span4Mux_v I__7870 (
            .O(N__33780),
            .I(N__33771));
    InMux I__7869 (
            .O(N__33779),
            .I(N__33766));
    InMux I__7868 (
            .O(N__33778),
            .I(N__33766));
    Span4Mux_h I__7867 (
            .O(N__33775),
            .I(N__33763));
    InMux I__7866 (
            .O(N__33774),
            .I(N__33760));
    Odrv4 I__7865 (
            .O(N__33771),
            .I(\this_ppu.N_510 ));
    LocalMux I__7864 (
            .O(N__33766),
            .I(\this_ppu.N_510 ));
    Odrv4 I__7863 (
            .O(N__33763),
            .I(\this_ppu.N_510 ));
    LocalMux I__7862 (
            .O(N__33760),
            .I(\this_ppu.N_510 ));
    InMux I__7861 (
            .O(N__33751),
            .I(N__33748));
    LocalMux I__7860 (
            .O(N__33748),
            .I(N__33742));
    InMux I__7859 (
            .O(N__33747),
            .I(N__33739));
    InMux I__7858 (
            .O(N__33746),
            .I(N__33734));
    InMux I__7857 (
            .O(N__33745),
            .I(N__33734));
    Span4Mux_h I__7856 (
            .O(N__33742),
            .I(N__33731));
    LocalMux I__7855 (
            .O(N__33739),
            .I(N__33726));
    LocalMux I__7854 (
            .O(N__33734),
            .I(N__33726));
    Sp12to4 I__7853 (
            .O(N__33731),
            .I(N__33721));
    Span12Mux_h I__7852 (
            .O(N__33726),
            .I(N__33721));
    Span12Mux_v I__7851 (
            .O(N__33721),
            .I(N__33718));
    Odrv12 I__7850 (
            .O(N__33718),
            .I(port_address_in_1));
    InMux I__7849 (
            .O(N__33715),
            .I(N__33710));
    InMux I__7848 (
            .O(N__33714),
            .I(N__33705));
    InMux I__7847 (
            .O(N__33713),
            .I(N__33705));
    LocalMux I__7846 (
            .O(N__33710),
            .I(\this_ppu.N_916 ));
    LocalMux I__7845 (
            .O(N__33705),
            .I(\this_ppu.N_916 ));
    InMux I__7844 (
            .O(N__33700),
            .I(N__33697));
    LocalMux I__7843 (
            .O(N__33697),
            .I(N__33694));
    Span4Mux_v I__7842 (
            .O(N__33694),
            .I(N__33691));
    Odrv4 I__7841 (
            .O(N__33691),
            .I(N_433));
    InMux I__7840 (
            .O(N__33688),
            .I(N__33685));
    LocalMux I__7839 (
            .O(N__33685),
            .I(N__33682));
    Span4Mux_v I__7838 (
            .O(N__33682),
            .I(N__33679));
    Span4Mux_h I__7837 (
            .O(N__33679),
            .I(N__33676));
    Odrv4 I__7836 (
            .O(N__33676),
            .I(N_438));
    InMux I__7835 (
            .O(N__33673),
            .I(N__33670));
    LocalMux I__7834 (
            .O(N__33670),
            .I(N__33667));
    Odrv12 I__7833 (
            .O(N__33667),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__7832 (
            .O(N__33664),
            .I(N__33661));
    LocalMux I__7831 (
            .O(N__33661),
            .I(N__33658));
    Odrv12 I__7830 (
            .O(N__33658),
            .I(M_this_oam_ram_write_data_12));
    CascadeMux I__7829 (
            .O(N__33655),
            .I(N__33652));
    InMux I__7828 (
            .O(N__33652),
            .I(N__33649));
    LocalMux I__7827 (
            .O(N__33649),
            .I(N__33646));
    Span4Mux_h I__7826 (
            .O(N__33646),
            .I(N__33643));
    Odrv4 I__7825 (
            .O(N__33643),
            .I(M_this_scroll_qZ0Z_2));
    CEMux I__7824 (
            .O(N__33640),
            .I(N__33637));
    LocalMux I__7823 (
            .O(N__33637),
            .I(N__33634));
    Span4Mux_v I__7822 (
            .O(N__33634),
            .I(N__33630));
    CEMux I__7821 (
            .O(N__33633),
            .I(N__33627));
    Span4Mux_h I__7820 (
            .O(N__33630),
            .I(N__33622));
    LocalMux I__7819 (
            .O(N__33627),
            .I(N__33622));
    Sp12to4 I__7818 (
            .O(N__33622),
            .I(N__33619));
    Odrv12 I__7817 (
            .O(N__33619),
            .I(N_1318_0));
    InMux I__7816 (
            .O(N__33616),
            .I(N__33613));
    LocalMux I__7815 (
            .O(N__33613),
            .I(M_this_data_tmp_qZ0Z_0));
    InMux I__7814 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__7813 (
            .O(N__33607),
            .I(N__33604));
    Span4Mux_h I__7812 (
            .O(N__33604),
            .I(N__33601));
    Odrv4 I__7811 (
            .O(N__33601),
            .I(M_this_oam_ram_write_data_0));
    InMux I__7810 (
            .O(N__33598),
            .I(N__33595));
    LocalMux I__7809 (
            .O(N__33595),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__7808 (
            .O(N__33592),
            .I(N__33589));
    LocalMux I__7807 (
            .O(N__33589),
            .I(N__33586));
    Span4Mux_h I__7806 (
            .O(N__33586),
            .I(N__33583));
    Odrv4 I__7805 (
            .O(N__33583),
            .I(M_this_oam_ram_write_data_1));
    InMux I__7804 (
            .O(N__33580),
            .I(N__33577));
    LocalMux I__7803 (
            .O(N__33577),
            .I(N__33574));
    Odrv12 I__7802 (
            .O(N__33574),
            .I(N_434));
    InMux I__7801 (
            .O(N__33571),
            .I(N__33568));
    LocalMux I__7800 (
            .O(N__33568),
            .I(N__33565));
    Odrv4 I__7799 (
            .O(N__33565),
            .I(\this_spr_ram.mem_out_bus5_3 ));
    InMux I__7798 (
            .O(N__33562),
            .I(N__33559));
    LocalMux I__7797 (
            .O(N__33559),
            .I(N__33556));
    Span4Mux_h I__7796 (
            .O(N__33556),
            .I(N__33553));
    Odrv4 I__7795 (
            .O(N__33553),
            .I(\this_spr_ram.mem_out_bus1_3 ));
    InMux I__7794 (
            .O(N__33550),
            .I(N__33547));
    LocalMux I__7793 (
            .O(N__33547),
            .I(N__33544));
    Span4Mux_h I__7792 (
            .O(N__33544),
            .I(N__33541));
    Odrv4 I__7791 (
            .O(N__33541),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ));
    CascadeMux I__7790 (
            .O(N__33538),
            .I(N__33534));
    CascadeMux I__7789 (
            .O(N__33537),
            .I(N__33531));
    InMux I__7788 (
            .O(N__33534),
            .I(N__33528));
    InMux I__7787 (
            .O(N__33531),
            .I(N__33524));
    LocalMux I__7786 (
            .O(N__33528),
            .I(N__33521));
    InMux I__7785 (
            .O(N__33527),
            .I(N__33518));
    LocalMux I__7784 (
            .O(N__33524),
            .I(\this_ppu.M_voffset_qZ0Z_2 ));
    Odrv12 I__7783 (
            .O(N__33521),
            .I(\this_ppu.M_voffset_qZ0Z_2 ));
    LocalMux I__7782 (
            .O(N__33518),
            .I(\this_ppu.M_voffset_qZ0Z_2 ));
    CascadeMux I__7781 (
            .O(N__33511),
            .I(N__33508));
    InMux I__7780 (
            .O(N__33508),
            .I(N__33505));
    LocalMux I__7779 (
            .O(N__33505),
            .I(\this_ppu.M_voffset_q_i_2 ));
    CascadeMux I__7778 (
            .O(N__33502),
            .I(N__33499));
    CascadeBuf I__7777 (
            .O(N__33499),
            .I(N__33496));
    CascadeMux I__7776 (
            .O(N__33496),
            .I(N__33493));
    InMux I__7775 (
            .O(N__33493),
            .I(N__33490));
    LocalMux I__7774 (
            .O(N__33490),
            .I(N__33486));
    CascadeMux I__7773 (
            .O(N__33489),
            .I(N__33483));
    Span4Mux_h I__7772 (
            .O(N__33486),
            .I(N__33480));
    InMux I__7771 (
            .O(N__33483),
            .I(N__33477));
    Span4Mux_h I__7770 (
            .O(N__33480),
            .I(N__33473));
    LocalMux I__7769 (
            .O(N__33477),
            .I(N__33470));
    InMux I__7768 (
            .O(N__33476),
            .I(N__33467));
    Span4Mux_h I__7767 (
            .O(N__33473),
            .I(N__33464));
    Odrv4 I__7766 (
            .O(N__33470),
            .I(M_this_ppu_map_addr_5));
    LocalMux I__7765 (
            .O(N__33467),
            .I(M_this_ppu_map_addr_5));
    Odrv4 I__7764 (
            .O(N__33464),
            .I(M_this_ppu_map_addr_5));
    CascadeMux I__7763 (
            .O(N__33457),
            .I(N__33454));
    InMux I__7762 (
            .O(N__33454),
            .I(N__33451));
    LocalMux I__7761 (
            .O(N__33451),
            .I(\this_ppu.M_this_ppu_map_addr_i_5 ));
    CascadeMux I__7760 (
            .O(N__33448),
            .I(N__33445));
    CascadeBuf I__7759 (
            .O(N__33445),
            .I(N__33442));
    CascadeMux I__7758 (
            .O(N__33442),
            .I(N__33439));
    InMux I__7757 (
            .O(N__33439),
            .I(N__33435));
    CascadeMux I__7756 (
            .O(N__33438),
            .I(N__33432));
    LocalMux I__7755 (
            .O(N__33435),
            .I(N__33429));
    InMux I__7754 (
            .O(N__33432),
            .I(N__33426));
    Span12Mux_s8_h I__7753 (
            .O(N__33429),
            .I(N__33422));
    LocalMux I__7752 (
            .O(N__33426),
            .I(N__33419));
    InMux I__7751 (
            .O(N__33425),
            .I(N__33416));
    Span12Mux_h I__7750 (
            .O(N__33422),
            .I(N__33413));
    Odrv12 I__7749 (
            .O(N__33419),
            .I(M_this_ppu_map_addr_6));
    LocalMux I__7748 (
            .O(N__33416),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__7747 (
            .O(N__33413),
            .I(M_this_ppu_map_addr_6));
    CascadeMux I__7746 (
            .O(N__33406),
            .I(N__33403));
    InMux I__7745 (
            .O(N__33403),
            .I(N__33400));
    LocalMux I__7744 (
            .O(N__33400),
            .I(\this_ppu.M_this_ppu_map_addr_i_6 ));
    CascadeMux I__7743 (
            .O(N__33397),
            .I(N__33394));
    CascadeBuf I__7742 (
            .O(N__33394),
            .I(N__33391));
    CascadeMux I__7741 (
            .O(N__33391),
            .I(N__33387));
    CascadeMux I__7740 (
            .O(N__33390),
            .I(N__33384));
    InMux I__7739 (
            .O(N__33387),
            .I(N__33381));
    InMux I__7738 (
            .O(N__33384),
            .I(N__33378));
    LocalMux I__7737 (
            .O(N__33381),
            .I(N__33374));
    LocalMux I__7736 (
            .O(N__33378),
            .I(N__33371));
    InMux I__7735 (
            .O(N__33377),
            .I(N__33368));
    Span12Mux_h I__7734 (
            .O(N__33374),
            .I(N__33365));
    Odrv4 I__7733 (
            .O(N__33371),
            .I(M_this_ppu_map_addr_7));
    LocalMux I__7732 (
            .O(N__33368),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__7731 (
            .O(N__33365),
            .I(M_this_ppu_map_addr_7));
    CascadeMux I__7730 (
            .O(N__33358),
            .I(N__33355));
    InMux I__7729 (
            .O(N__33355),
            .I(N__33352));
    LocalMux I__7728 (
            .O(N__33352),
            .I(\this_ppu.M_this_ppu_map_addr_i_7 ));
    CascadeMux I__7727 (
            .O(N__33349),
            .I(N__33346));
    CascadeBuf I__7726 (
            .O(N__33346),
            .I(N__33342));
    CascadeMux I__7725 (
            .O(N__33345),
            .I(N__33339));
    CascadeMux I__7724 (
            .O(N__33342),
            .I(N__33336));
    InMux I__7723 (
            .O(N__33339),
            .I(N__33333));
    InMux I__7722 (
            .O(N__33336),
            .I(N__33330));
    LocalMux I__7721 (
            .O(N__33333),
            .I(N__33327));
    LocalMux I__7720 (
            .O(N__33330),
            .I(N__33323));
    Span4Mux_h I__7719 (
            .O(N__33327),
            .I(N__33320));
    InMux I__7718 (
            .O(N__33326),
            .I(N__33317));
    Span12Mux_s10_h I__7717 (
            .O(N__33323),
            .I(N__33314));
    Odrv4 I__7716 (
            .O(N__33320),
            .I(M_this_ppu_map_addr_8));
    LocalMux I__7715 (
            .O(N__33317),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__7714 (
            .O(N__33314),
            .I(M_this_ppu_map_addr_8));
    CascadeMux I__7713 (
            .O(N__33307),
            .I(N__33304));
    InMux I__7712 (
            .O(N__33304),
            .I(N__33301));
    LocalMux I__7711 (
            .O(N__33301),
            .I(\this_ppu.M_this_ppu_map_addr_i_8 ));
    CascadeMux I__7710 (
            .O(N__33298),
            .I(N__33295));
    CascadeBuf I__7709 (
            .O(N__33295),
            .I(N__33292));
    CascadeMux I__7708 (
            .O(N__33292),
            .I(N__33288));
    CascadeMux I__7707 (
            .O(N__33291),
            .I(N__33285));
    InMux I__7706 (
            .O(N__33288),
            .I(N__33282));
    InMux I__7705 (
            .O(N__33285),
            .I(N__33279));
    LocalMux I__7704 (
            .O(N__33282),
            .I(N__33275));
    LocalMux I__7703 (
            .O(N__33279),
            .I(N__33272));
    InMux I__7702 (
            .O(N__33278),
            .I(N__33269));
    Span12Mux_s9_h I__7701 (
            .O(N__33275),
            .I(N__33266));
    Odrv12 I__7700 (
            .O(N__33272),
            .I(M_this_ppu_map_addr_9));
    LocalMux I__7699 (
            .O(N__33269),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__7698 (
            .O(N__33266),
            .I(M_this_ppu_map_addr_9));
    CascadeMux I__7697 (
            .O(N__33259),
            .I(N__33256));
    InMux I__7696 (
            .O(N__33256),
            .I(N__33253));
    LocalMux I__7695 (
            .O(N__33253),
            .I(\this_ppu.M_this_ppu_map_addr_i_9 ));
    CascadeMux I__7694 (
            .O(N__33250),
            .I(N__33247));
    InMux I__7693 (
            .O(N__33247),
            .I(N__33244));
    LocalMux I__7692 (
            .O(N__33244),
            .I(N__33240));
    InMux I__7691 (
            .O(N__33243),
            .I(N__33237));
    Odrv4 I__7690 (
            .O(N__33240),
            .I(\this_ppu.M_voffset_qZ0Z_8 ));
    LocalMux I__7689 (
            .O(N__33237),
            .I(\this_ppu.M_voffset_qZ0Z_8 ));
    InMux I__7688 (
            .O(N__33232),
            .I(N__33229));
    LocalMux I__7687 (
            .O(N__33229),
            .I(\this_ppu.M_voffset_q_i_8 ));
    InMux I__7686 (
            .O(N__33226),
            .I(\this_ppu.un1_M_voffset_q_cry_8 ));
    InMux I__7685 (
            .O(N__33223),
            .I(N__33220));
    LocalMux I__7684 (
            .O(N__33220),
            .I(N__33217));
    Span4Mux_v I__7683 (
            .O(N__33217),
            .I(N__33212));
    InMux I__7682 (
            .O(N__33216),
            .I(N__33209));
    InMux I__7681 (
            .O(N__33215),
            .I(N__33206));
    Span4Mux_v I__7680 (
            .O(N__33212),
            .I(N__33203));
    LocalMux I__7679 (
            .O(N__33209),
            .I(N__33198));
    LocalMux I__7678 (
            .O(N__33206),
            .I(N__33198));
    Span4Mux_v I__7677 (
            .O(N__33203),
            .I(N__33195));
    Span4Mux_h I__7676 (
            .O(N__33198),
            .I(N__33192));
    Odrv4 I__7675 (
            .O(N__33195),
            .I(\this_ppu.M_state_d14_1 ));
    Odrv4 I__7674 (
            .O(N__33192),
            .I(\this_ppu.M_state_d14_1 ));
    CascadeMux I__7673 (
            .O(N__33187),
            .I(N__33184));
    InMux I__7672 (
            .O(N__33184),
            .I(N__33181));
    LocalMux I__7671 (
            .O(N__33181),
            .I(N__33177));
    CascadeMux I__7670 (
            .O(N__33180),
            .I(N__33174));
    Span4Mux_v I__7669 (
            .O(N__33177),
            .I(N__33171));
    InMux I__7668 (
            .O(N__33174),
            .I(N__33168));
    Odrv4 I__7667 (
            .O(N__33171),
            .I(M_this_scroll_qZ0Z_0));
    LocalMux I__7666 (
            .O(N__33168),
            .I(M_this_scroll_qZ0Z_0));
    CascadeMux I__7665 (
            .O(N__33163),
            .I(N__33160));
    InMux I__7664 (
            .O(N__33160),
            .I(N__33157));
    LocalMux I__7663 (
            .O(N__33157),
            .I(M_this_scroll_qZ0Z_1));
    CascadeMux I__7662 (
            .O(N__33154),
            .I(N__33151));
    InMux I__7661 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__7660 (
            .O(N__33148),
            .I(M_this_scroll_qZ0Z_5));
    CascadeMux I__7659 (
            .O(N__33145),
            .I(N__33142));
    InMux I__7658 (
            .O(N__33142),
            .I(N__33139));
    LocalMux I__7657 (
            .O(N__33139),
            .I(M_this_scroll_qZ0Z_3));
    InMux I__7656 (
            .O(N__33136),
            .I(N__33133));
    LocalMux I__7655 (
            .O(N__33133),
            .I(M_this_scroll_qZ0Z_4));
    InMux I__7654 (
            .O(N__33130),
            .I(N__33127));
    LocalMux I__7653 (
            .O(N__33127),
            .I(M_this_scroll_qZ0Z_6));
    CascadeMux I__7652 (
            .O(N__33124),
            .I(N__33121));
    InMux I__7651 (
            .O(N__33121),
            .I(N__33118));
    LocalMux I__7650 (
            .O(N__33118),
            .I(M_this_scroll_qZ0Z_7));
    CascadeMux I__7649 (
            .O(N__33115),
            .I(N__33112));
    InMux I__7648 (
            .O(N__33112),
            .I(N__33109));
    LocalMux I__7647 (
            .O(N__33109),
            .I(\this_ppu.M_voffset_q_i_0 ));
    CascadeMux I__7646 (
            .O(N__33106),
            .I(N__33103));
    InMux I__7645 (
            .O(N__33103),
            .I(N__33099));
    InMux I__7644 (
            .O(N__33102),
            .I(N__33095));
    LocalMux I__7643 (
            .O(N__33099),
            .I(N__33092));
    InMux I__7642 (
            .O(N__33098),
            .I(N__33089));
    LocalMux I__7641 (
            .O(N__33095),
            .I(\this_ppu.M_voffset_qZ0Z_1 ));
    Odrv12 I__7640 (
            .O(N__33092),
            .I(\this_ppu.M_voffset_qZ0Z_1 ));
    LocalMux I__7639 (
            .O(N__33089),
            .I(\this_ppu.M_voffset_qZ0Z_1 ));
    CascadeMux I__7638 (
            .O(N__33082),
            .I(N__33079));
    InMux I__7637 (
            .O(N__33079),
            .I(N__33076));
    LocalMux I__7636 (
            .O(N__33076),
            .I(\this_ppu.M_voffset_q_i_1 ));
    CascadeMux I__7635 (
            .O(N__33073),
            .I(N__33070));
    CascadeBuf I__7634 (
            .O(N__33070),
            .I(N__33067));
    CascadeMux I__7633 (
            .O(N__33067),
            .I(N__33064));
    InMux I__7632 (
            .O(N__33064),
            .I(N__33060));
    CascadeMux I__7631 (
            .O(N__33063),
            .I(N__33057));
    LocalMux I__7630 (
            .O(N__33060),
            .I(N__33054));
    InMux I__7629 (
            .O(N__33057),
            .I(N__33051));
    Span4Mux_v I__7628 (
            .O(N__33054),
            .I(N__33046));
    LocalMux I__7627 (
            .O(N__33051),
            .I(N__33043));
    InMux I__7626 (
            .O(N__33050),
            .I(N__33040));
    CascadeMux I__7625 (
            .O(N__33049),
            .I(N__33037));
    Span4Mux_h I__7624 (
            .O(N__33046),
            .I(N__33034));
    Span4Mux_v I__7623 (
            .O(N__33043),
            .I(N__33029));
    LocalMux I__7622 (
            .O(N__33040),
            .I(N__33029));
    InMux I__7621 (
            .O(N__33037),
            .I(N__33026));
    Span4Mux_h I__7620 (
            .O(N__33034),
            .I(N__33023));
    Span4Mux_h I__7619 (
            .O(N__33029),
            .I(N__33020));
    LocalMux I__7618 (
            .O(N__33026),
            .I(N__33015));
    Span4Mux_h I__7617 (
            .O(N__33023),
            .I(N__33015));
    Odrv4 I__7616 (
            .O(N__33020),
            .I(M_this_ppu_map_addr_0));
    Odrv4 I__7615 (
            .O(N__33015),
            .I(M_this_ppu_map_addr_0));
    InMux I__7614 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__7613 (
            .O(N__33007),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0 ));
    CascadeMux I__7612 (
            .O(N__33004),
            .I(N__33001));
    CascadeBuf I__7611 (
            .O(N__33001),
            .I(N__32998));
    CascadeMux I__7610 (
            .O(N__32998),
            .I(N__32995));
    InMux I__7609 (
            .O(N__32995),
            .I(N__32991));
    CascadeMux I__7608 (
            .O(N__32994),
            .I(N__32986));
    LocalMux I__7607 (
            .O(N__32991),
            .I(N__32982));
    InMux I__7606 (
            .O(N__32990),
            .I(N__32979));
    InMux I__7605 (
            .O(N__32989),
            .I(N__32975));
    InMux I__7604 (
            .O(N__32986),
            .I(N__32972));
    InMux I__7603 (
            .O(N__32985),
            .I(N__32969));
    Span4Mux_h I__7602 (
            .O(N__32982),
            .I(N__32966));
    LocalMux I__7601 (
            .O(N__32979),
            .I(N__32963));
    InMux I__7600 (
            .O(N__32978),
            .I(N__32960));
    LocalMux I__7599 (
            .O(N__32975),
            .I(N__32955));
    LocalMux I__7598 (
            .O(N__32972),
            .I(N__32955));
    LocalMux I__7597 (
            .O(N__32969),
            .I(N__32952));
    Sp12to4 I__7596 (
            .O(N__32966),
            .I(N__32949));
    Span4Mux_h I__7595 (
            .O(N__32963),
            .I(N__32946));
    LocalMux I__7594 (
            .O(N__32960),
            .I(N__32943));
    Span4Mux_v I__7593 (
            .O(N__32955),
            .I(N__32940));
    Span4Mux_v I__7592 (
            .O(N__32952),
            .I(N__32937));
    Span12Mux_v I__7591 (
            .O(N__32949),
            .I(N__32934));
    Odrv4 I__7590 (
            .O(N__32946),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__7589 (
            .O(N__32943),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__7588 (
            .O(N__32940),
            .I(M_this_ppu_map_addr_1));
    Odrv4 I__7587 (
            .O(N__32937),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__7586 (
            .O(N__32934),
            .I(M_this_ppu_map_addr_1));
    CascadeMux I__7585 (
            .O(N__32923),
            .I(N__32920));
    CascadeBuf I__7584 (
            .O(N__32920),
            .I(N__32916));
    InMux I__7583 (
            .O(N__32919),
            .I(N__32912));
    CascadeMux I__7582 (
            .O(N__32916),
            .I(N__32909));
    CascadeMux I__7581 (
            .O(N__32915),
            .I(N__32906));
    LocalMux I__7580 (
            .O(N__32912),
            .I(N__32903));
    InMux I__7579 (
            .O(N__32909),
            .I(N__32899));
    InMux I__7578 (
            .O(N__32906),
            .I(N__32896));
    Span4Mux_v I__7577 (
            .O(N__32903),
            .I(N__32893));
    InMux I__7576 (
            .O(N__32902),
            .I(N__32890));
    LocalMux I__7575 (
            .O(N__32899),
            .I(N__32887));
    LocalMux I__7574 (
            .O(N__32896),
            .I(N__32884));
    Span4Mux_h I__7573 (
            .O(N__32893),
            .I(N__32879));
    LocalMux I__7572 (
            .O(N__32890),
            .I(N__32879));
    Sp12to4 I__7571 (
            .O(N__32887),
            .I(N__32876));
    Span4Mux_h I__7570 (
            .O(N__32884),
            .I(N__32873));
    Span4Mux_h I__7569 (
            .O(N__32879),
            .I(N__32870));
    Span12Mux_h I__7568 (
            .O(N__32876),
            .I(N__32867));
    Odrv4 I__7567 (
            .O(N__32873),
            .I(M_this_ppu_map_addr_3));
    Odrv4 I__7566 (
            .O(N__32870),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__7565 (
            .O(N__32867),
            .I(M_this_ppu_map_addr_3));
    InMux I__7564 (
            .O(N__32860),
            .I(N__32857));
    LocalMux I__7563 (
            .O(N__32857),
            .I(N__32853));
    CascadeMux I__7562 (
            .O(N__32856),
            .I(N__32850));
    Span4Mux_h I__7561 (
            .O(N__32853),
            .I(N__32847));
    InMux I__7560 (
            .O(N__32850),
            .I(N__32844));
    Odrv4 I__7559 (
            .O(N__32847),
            .I(\this_ppu.read_data_RNI3DGK1_14 ));
    LocalMux I__7558 (
            .O(N__32844),
            .I(\this_ppu.read_data_RNI3DGK1_14 ));
    InMux I__7557 (
            .O(N__32839),
            .I(N__32836));
    LocalMux I__7556 (
            .O(N__32836),
            .I(N__32833));
    Odrv4 I__7555 (
            .O(N__32833),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0 ));
    CascadeMux I__7554 (
            .O(N__32830),
            .I(N__32827));
    InMux I__7553 (
            .O(N__32827),
            .I(N__32823));
    InMux I__7552 (
            .O(N__32826),
            .I(N__32819));
    LocalMux I__7551 (
            .O(N__32823),
            .I(N__32816));
    InMux I__7550 (
            .O(N__32822),
            .I(N__32813));
    LocalMux I__7549 (
            .O(N__32819),
            .I(N__32806));
    Span4Mux_v I__7548 (
            .O(N__32816),
            .I(N__32806));
    LocalMux I__7547 (
            .O(N__32813),
            .I(N__32806));
    Span4Mux_h I__7546 (
            .O(N__32806),
            .I(N__32803));
    Odrv4 I__7545 (
            .O(N__32803),
            .I(\this_ppu.M_hoffset_qZ0Z_8 ));
    InMux I__7544 (
            .O(N__32800),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_8 ));
    CascadeMux I__7543 (
            .O(N__32797),
            .I(N__32794));
    InMux I__7542 (
            .O(N__32794),
            .I(N__32791));
    LocalMux I__7541 (
            .O(N__32791),
            .I(N__32788));
    Span4Mux_h I__7540 (
            .O(N__32788),
            .I(N__32785));
    Odrv4 I__7539 (
            .O(N__32785),
            .I(\this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO ));
    InMux I__7538 (
            .O(N__32782),
            .I(N__32779));
    LocalMux I__7537 (
            .O(N__32779),
            .I(N__32776));
    Span4Mux_h I__7536 (
            .O(N__32776),
            .I(N__32773));
    Odrv4 I__7535 (
            .O(N__32773),
            .I(\this_ppu.oam_cache.mem_18 ));
    InMux I__7534 (
            .O(N__32770),
            .I(N__32767));
    LocalMux I__7533 (
            .O(N__32767),
            .I(\this_ppu.M_oam_cache_read_data_18 ));
    InMux I__7532 (
            .O(N__32764),
            .I(N__32761));
    LocalMux I__7531 (
            .O(N__32761),
            .I(\this_ppu.un1_oam_data_1_6 ));
    InMux I__7530 (
            .O(N__32758),
            .I(N__32755));
    LocalMux I__7529 (
            .O(N__32755),
            .I(\this_ppu.un1_oam_data_1_8 ));
    InMux I__7528 (
            .O(N__32752),
            .I(N__32749));
    LocalMux I__7527 (
            .O(N__32749),
            .I(\this_ppu.un1_oam_data_1_7 ));
    InMux I__7526 (
            .O(N__32746),
            .I(N__32743));
    LocalMux I__7525 (
            .O(N__32743),
            .I(\this_ppu.un1_oam_data_1_5 ));
    CascadeMux I__7524 (
            .O(N__32740),
            .I(N__32736));
    CascadeMux I__7523 (
            .O(N__32739),
            .I(N__32733));
    InMux I__7522 (
            .O(N__32736),
            .I(N__32730));
    InMux I__7521 (
            .O(N__32733),
            .I(N__32727));
    LocalMux I__7520 (
            .O(N__32730),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    LocalMux I__7519 (
            .O(N__32727),
            .I(\this_ppu.M_this_ppu_map_addr_i_2 ));
    CascadeMux I__7518 (
            .O(N__32722),
            .I(N__32718));
    CascadeMux I__7517 (
            .O(N__32721),
            .I(N__32715));
    InMux I__7516 (
            .O(N__32718),
            .I(N__32712));
    InMux I__7515 (
            .O(N__32715),
            .I(N__32709));
    LocalMux I__7514 (
            .O(N__32712),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    LocalMux I__7513 (
            .O(N__32709),
            .I(\this_ppu.M_this_ppu_map_addr_i_3 ));
    InMux I__7512 (
            .O(N__32704),
            .I(N__32700));
    InMux I__7511 (
            .O(N__32703),
            .I(N__32697));
    LocalMux I__7510 (
            .O(N__32700),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    LocalMux I__7509 (
            .O(N__32697),
            .I(\this_ppu.M_this_ppu_map_addr_i_4 ));
    InMux I__7508 (
            .O(N__32692),
            .I(bfn_22_19_0_));
    InMux I__7507 (
            .O(N__32689),
            .I(N__32686));
    LocalMux I__7506 (
            .O(N__32686),
            .I(N__32683));
    Span4Mux_h I__7505 (
            .O(N__32683),
            .I(N__32680));
    Odrv4 I__7504 (
            .O(N__32680),
            .I(\this_ppu.vspr16_0 ));
    InMux I__7503 (
            .O(N__32677),
            .I(N__32674));
    LocalMux I__7502 (
            .O(N__32674),
            .I(N__32671));
    Span4Mux_h I__7501 (
            .O(N__32671),
            .I(N__32668));
    Odrv4 I__7500 (
            .O(N__32668),
            .I(\this_ppu.un1_M_oam_cache_read_data_ac0_13_i ));
    CascadeMux I__7499 (
            .O(N__32665),
            .I(N__32662));
    InMux I__7498 (
            .O(N__32662),
            .I(N__32659));
    LocalMux I__7497 (
            .O(N__32659),
            .I(N__32656));
    Odrv4 I__7496 (
            .O(N__32656),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0 ));
    CascadeMux I__7495 (
            .O(N__32653),
            .I(N__32650));
    InMux I__7494 (
            .O(N__32650),
            .I(N__32647));
    LocalMux I__7493 (
            .O(N__32647),
            .I(N__32644));
    Odrv12 I__7492 (
            .O(N__32644),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0 ));
    CascadeMux I__7491 (
            .O(N__32641),
            .I(N__32638));
    InMux I__7490 (
            .O(N__32638),
            .I(N__32635));
    LocalMux I__7489 (
            .O(N__32635),
            .I(N__32632));
    Odrv4 I__7488 (
            .O(N__32632),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0 ));
    CascadeMux I__7487 (
            .O(N__32629),
            .I(N__32622));
    InMux I__7486 (
            .O(N__32628),
            .I(N__32617));
    InMux I__7485 (
            .O(N__32627),
            .I(N__32617));
    InMux I__7484 (
            .O(N__32626),
            .I(N__32614));
    InMux I__7483 (
            .O(N__32625),
            .I(N__32609));
    InMux I__7482 (
            .O(N__32622),
            .I(N__32609));
    LocalMux I__7481 (
            .O(N__32617),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__7480 (
            .O(N__32614),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__7479 (
            .O(N__32609),
            .I(M_this_state_qZ0Z_3));
    InMux I__7478 (
            .O(N__32602),
            .I(N__32598));
    CascadeMux I__7477 (
            .O(N__32601),
            .I(N__32594));
    LocalMux I__7476 (
            .O(N__32598),
            .I(N__32591));
    CascadeMux I__7475 (
            .O(N__32597),
            .I(N__32587));
    InMux I__7474 (
            .O(N__32594),
            .I(N__32583));
    Span4Mux_v I__7473 (
            .O(N__32591),
            .I(N__32580));
    InMux I__7472 (
            .O(N__32590),
            .I(N__32575));
    InMux I__7471 (
            .O(N__32587),
            .I(N__32575));
    InMux I__7470 (
            .O(N__32586),
            .I(N__32572));
    LocalMux I__7469 (
            .O(N__32583),
            .I(M_this_state_qZ0Z_2));
    Odrv4 I__7468 (
            .O(N__32580),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__7467 (
            .O(N__32575),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__7466 (
            .O(N__32572),
            .I(M_this_state_qZ0Z_2));
    InMux I__7465 (
            .O(N__32563),
            .I(N__32560));
    LocalMux I__7464 (
            .O(N__32560),
            .I(\this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0 ));
    CascadeMux I__7463 (
            .O(N__32557),
            .I(\this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_ ));
    InMux I__7462 (
            .O(N__32554),
            .I(N__32551));
    LocalMux I__7461 (
            .O(N__32551),
            .I(\this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0 ));
    InMux I__7460 (
            .O(N__32548),
            .I(N__32545));
    LocalMux I__7459 (
            .O(N__32545),
            .I(N__32542));
    Odrv4 I__7458 (
            .O(N__32542),
            .I(\this_ppu.N_416 ));
    CascadeMux I__7457 (
            .O(N__32539),
            .I(N__32535));
    CascadeMux I__7456 (
            .O(N__32538),
            .I(N__32532));
    InMux I__7455 (
            .O(N__32535),
            .I(N__32529));
    InMux I__7454 (
            .O(N__32532),
            .I(N__32526));
    LocalMux I__7453 (
            .O(N__32529),
            .I(\this_ppu.M_hoffset_q_i_0 ));
    LocalMux I__7452 (
            .O(N__32526),
            .I(\this_ppu.M_hoffset_q_i_0 ));
    CascadeMux I__7451 (
            .O(N__32521),
            .I(N__32517));
    CascadeMux I__7450 (
            .O(N__32520),
            .I(N__32514));
    InMux I__7449 (
            .O(N__32517),
            .I(N__32511));
    InMux I__7448 (
            .O(N__32514),
            .I(N__32508));
    LocalMux I__7447 (
            .O(N__32511),
            .I(\this_ppu.M_hoffset_q_i_1 ));
    LocalMux I__7446 (
            .O(N__32508),
            .I(\this_ppu.M_hoffset_q_i_1 ));
    CascadeMux I__7445 (
            .O(N__32503),
            .I(N__32499));
    CascadeMux I__7444 (
            .O(N__32502),
            .I(N__32496));
    InMux I__7443 (
            .O(N__32499),
            .I(N__32493));
    InMux I__7442 (
            .O(N__32496),
            .I(N__32490));
    LocalMux I__7441 (
            .O(N__32493),
            .I(\this_ppu.M_hoffset_q_i_2 ));
    LocalMux I__7440 (
            .O(N__32490),
            .I(\this_ppu.M_hoffset_q_i_2 ));
    CascadeMux I__7439 (
            .O(N__32485),
            .I(N__32482));
    InMux I__7438 (
            .O(N__32482),
            .I(N__32478));
    CascadeMux I__7437 (
            .O(N__32481),
            .I(N__32475));
    LocalMux I__7436 (
            .O(N__32478),
            .I(N__32472));
    InMux I__7435 (
            .O(N__32475),
            .I(N__32469));
    Odrv4 I__7434 (
            .O(N__32472),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    LocalMux I__7433 (
            .O(N__32469),
            .I(\this_ppu.M_this_ppu_map_addr_i_0 ));
    CascadeMux I__7432 (
            .O(N__32464),
            .I(N__32460));
    CascadeMux I__7431 (
            .O(N__32463),
            .I(N__32457));
    InMux I__7430 (
            .O(N__32460),
            .I(N__32454));
    InMux I__7429 (
            .O(N__32457),
            .I(N__32451));
    LocalMux I__7428 (
            .O(N__32454),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    LocalMux I__7427 (
            .O(N__32451),
            .I(\this_ppu.M_this_ppu_map_addr_i_1 ));
    CEMux I__7426 (
            .O(N__32446),
            .I(N__32443));
    LocalMux I__7425 (
            .O(N__32443),
            .I(N__32439));
    CEMux I__7424 (
            .O(N__32442),
            .I(N__32434));
    Span4Mux_v I__7423 (
            .O(N__32439),
            .I(N__32431));
    CEMux I__7422 (
            .O(N__32438),
            .I(N__32428));
    CEMux I__7421 (
            .O(N__32437),
            .I(N__32424));
    LocalMux I__7420 (
            .O(N__32434),
            .I(N__32419));
    Span4Mux_h I__7419 (
            .O(N__32431),
            .I(N__32414));
    LocalMux I__7418 (
            .O(N__32428),
            .I(N__32414));
    CEMux I__7417 (
            .O(N__32427),
            .I(N__32411));
    LocalMux I__7416 (
            .O(N__32424),
            .I(N__32408));
    CEMux I__7415 (
            .O(N__32423),
            .I(N__32405));
    CEMux I__7414 (
            .O(N__32422),
            .I(N__32402));
    Span4Mux_h I__7413 (
            .O(N__32419),
            .I(N__32395));
    Span4Mux_v I__7412 (
            .O(N__32414),
            .I(N__32395));
    LocalMux I__7411 (
            .O(N__32411),
            .I(N__32395));
    Span4Mux_v I__7410 (
            .O(N__32408),
            .I(N__32390));
    LocalMux I__7409 (
            .O(N__32405),
            .I(N__32390));
    LocalMux I__7408 (
            .O(N__32402),
            .I(N__32387));
    Span4Mux_h I__7407 (
            .O(N__32395),
            .I(N__32384));
    Span4Mux_h I__7406 (
            .O(N__32390),
            .I(N__32381));
    Span4Mux_v I__7405 (
            .O(N__32387),
            .I(N__32378));
    Span4Mux_v I__7404 (
            .O(N__32384),
            .I(N__32375));
    Span4Mux_v I__7403 (
            .O(N__32381),
            .I(N__32370));
    Span4Mux_h I__7402 (
            .O(N__32378),
            .I(N__32370));
    Odrv4 I__7401 (
            .O(N__32375),
            .I(N_1286_0));
    Odrv4 I__7400 (
            .O(N__32370),
            .I(N_1286_0));
    InMux I__7399 (
            .O(N__32365),
            .I(N__32362));
    LocalMux I__7398 (
            .O(N__32362),
            .I(N__32359));
    Span12Mux_h I__7397 (
            .O(N__32359),
            .I(N__32356));
    Span12Mux_v I__7396 (
            .O(N__32356),
            .I(N__32353));
    Odrv12 I__7395 (
            .O(N__32353),
            .I(M_this_map_ram_read_data_7));
    CascadeMux I__7394 (
            .O(N__32350),
            .I(N__32347));
    InMux I__7393 (
            .O(N__32347),
            .I(N__32343));
    CascadeMux I__7392 (
            .O(N__32346),
            .I(N__32340));
    LocalMux I__7391 (
            .O(N__32343),
            .I(N__32337));
    InMux I__7390 (
            .O(N__32340),
            .I(N__32334));
    Span4Mux_v I__7389 (
            .O(N__32337),
            .I(N__32331));
    LocalMux I__7388 (
            .O(N__32334),
            .I(N__32328));
    Span4Mux_v I__7387 (
            .O(N__32331),
            .I(N__32325));
    Span4Mux_v I__7386 (
            .O(N__32328),
            .I(N__32322));
    Odrv4 I__7385 (
            .O(N__32325),
            .I(\this_ppu.N_511 ));
    Odrv4 I__7384 (
            .O(N__32322),
            .I(\this_ppu.N_511 ));
    CascadeMux I__7383 (
            .O(N__32317),
            .I(\this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_ ));
    InMux I__7382 (
            .O(N__32314),
            .I(N__32311));
    LocalMux I__7381 (
            .O(N__32311),
            .I(N__32306));
    InMux I__7380 (
            .O(N__32310),
            .I(N__32303));
    InMux I__7379 (
            .O(N__32309),
            .I(N__32298));
    Span4Mux_h I__7378 (
            .O(N__32306),
            .I(N__32295));
    LocalMux I__7377 (
            .O(N__32303),
            .I(N__32292));
    InMux I__7376 (
            .O(N__32302),
            .I(N__32289));
    InMux I__7375 (
            .O(N__32301),
            .I(N__32286));
    LocalMux I__7374 (
            .O(N__32298),
            .I(M_this_state_qZ0Z_6));
    Odrv4 I__7373 (
            .O(N__32295),
            .I(M_this_state_qZ0Z_6));
    Odrv12 I__7372 (
            .O(N__32292),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__7371 (
            .O(N__32289),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__7370 (
            .O(N__32286),
            .I(M_this_state_qZ0Z_6));
    CascadeMux I__7369 (
            .O(N__32275),
            .I(N__32272));
    InMux I__7368 (
            .O(N__32272),
            .I(N__32269));
    LocalMux I__7367 (
            .O(N__32269),
            .I(N__32263));
    InMux I__7366 (
            .O(N__32268),
            .I(N__32257));
    InMux I__7365 (
            .O(N__32267),
            .I(N__32252));
    InMux I__7364 (
            .O(N__32266),
            .I(N__32252));
    Span4Mux_h I__7363 (
            .O(N__32263),
            .I(N__32249));
    InMux I__7362 (
            .O(N__32262),
            .I(N__32246));
    InMux I__7361 (
            .O(N__32261),
            .I(N__32241));
    InMux I__7360 (
            .O(N__32260),
            .I(N__32241));
    LocalMux I__7359 (
            .O(N__32257),
            .I(N__32238));
    LocalMux I__7358 (
            .O(N__32252),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__7357 (
            .O(N__32249),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__7356 (
            .O(N__32246),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__7355 (
            .O(N__32241),
            .I(M_this_state_qZ0Z_7));
    Odrv4 I__7354 (
            .O(N__32238),
            .I(M_this_state_qZ0Z_7));
    InMux I__7353 (
            .O(N__32227),
            .I(N__32224));
    LocalMux I__7352 (
            .O(N__32224),
            .I(this_ppu_un20_i_a4_0_a3_0_a2_1_1));
    InMux I__7351 (
            .O(N__32221),
            .I(N__32218));
    LocalMux I__7350 (
            .O(N__32218),
            .I(N__32214));
    InMux I__7349 (
            .O(N__32217),
            .I(N__32211));
    Span12Mux_v I__7348 (
            .O(N__32214),
            .I(N__32208));
    LocalMux I__7347 (
            .O(N__32211),
            .I(N__32205));
    Span12Mux_h I__7346 (
            .O(N__32208),
            .I(N__32202));
    Span4Mux_v I__7345 (
            .O(N__32205),
            .I(N__32199));
    Odrv12 I__7344 (
            .O(N__32202),
            .I(port_rw_in));
    Odrv4 I__7343 (
            .O(N__32199),
            .I(port_rw_in));
    CascadeMux I__7342 (
            .O(N__32194),
            .I(N__32190));
    InMux I__7341 (
            .O(N__32193),
            .I(N__32186));
    InMux I__7340 (
            .O(N__32190),
            .I(N__32180));
    CascadeMux I__7339 (
            .O(N__32189),
            .I(N__32177));
    LocalMux I__7338 (
            .O(N__32186),
            .I(N__32174));
    InMux I__7337 (
            .O(N__32185),
            .I(N__32171));
    InMux I__7336 (
            .O(N__32184),
            .I(N__32168));
    InMux I__7335 (
            .O(N__32183),
            .I(N__32165));
    LocalMux I__7334 (
            .O(N__32180),
            .I(N__32162));
    InMux I__7333 (
            .O(N__32177),
            .I(N__32159));
    Span4Mux_v I__7332 (
            .O(N__32174),
            .I(N__32152));
    LocalMux I__7331 (
            .O(N__32171),
            .I(N__32152));
    LocalMux I__7330 (
            .O(N__32168),
            .I(N__32152));
    LocalMux I__7329 (
            .O(N__32165),
            .I(N__32149));
    Span4Mux_v I__7328 (
            .O(N__32162),
            .I(N__32142));
    LocalMux I__7327 (
            .O(N__32159),
            .I(N__32142));
    Span4Mux_h I__7326 (
            .O(N__32152),
            .I(N__32142));
    Odrv4 I__7325 (
            .O(N__32149),
            .I(\this_ppu.N_321_0 ));
    Odrv4 I__7324 (
            .O(N__32142),
            .I(\this_ppu.N_321_0 ));
    CascadeMux I__7323 (
            .O(N__32137),
            .I(N__32133));
    InMux I__7322 (
            .O(N__32136),
            .I(N__32129));
    InMux I__7321 (
            .O(N__32133),
            .I(N__32124));
    InMux I__7320 (
            .O(N__32132),
            .I(N__32124));
    LocalMux I__7319 (
            .O(N__32129),
            .I(N__32118));
    LocalMux I__7318 (
            .O(N__32124),
            .I(N__32115));
    InMux I__7317 (
            .O(N__32123),
            .I(N__32112));
    CascadeMux I__7316 (
            .O(N__32122),
            .I(N__32108));
    InMux I__7315 (
            .O(N__32121),
            .I(N__32104));
    Span4Mux_h I__7314 (
            .O(N__32118),
            .I(N__32097));
    Span4Mux_v I__7313 (
            .O(N__32115),
            .I(N__32097));
    LocalMux I__7312 (
            .O(N__32112),
            .I(N__32097));
    InMux I__7311 (
            .O(N__32111),
            .I(N__32094));
    InMux I__7310 (
            .O(N__32108),
            .I(N__32089));
    InMux I__7309 (
            .O(N__32107),
            .I(N__32089));
    LocalMux I__7308 (
            .O(N__32104),
            .I(\this_ppu.N_328_0 ));
    Odrv4 I__7307 (
            .O(N__32097),
            .I(\this_ppu.N_328_0 ));
    LocalMux I__7306 (
            .O(N__32094),
            .I(\this_ppu.N_328_0 ));
    LocalMux I__7305 (
            .O(N__32089),
            .I(\this_ppu.N_328_0 ));
    InMux I__7304 (
            .O(N__32080),
            .I(\this_ppu.un1_M_voffset_d_cry_5 ));
    InMux I__7303 (
            .O(N__32077),
            .I(N__32073));
    InMux I__7302 (
            .O(N__32076),
            .I(N__32070));
    LocalMux I__7301 (
            .O(N__32073),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    LocalMux I__7300 (
            .O(N__32070),
            .I(\this_ppu.M_vaddress_qZ0Z_7 ));
    InMux I__7299 (
            .O(N__32065),
            .I(\this_ppu.un1_M_voffset_d_cry_6 ));
    InMux I__7298 (
            .O(N__32062),
            .I(bfn_21_24_0_));
    CEMux I__7297 (
            .O(N__32059),
            .I(N__32054));
    CEMux I__7296 (
            .O(N__32058),
            .I(N__32051));
    CEMux I__7295 (
            .O(N__32057),
            .I(N__32047));
    LocalMux I__7294 (
            .O(N__32054),
            .I(N__32044));
    LocalMux I__7293 (
            .O(N__32051),
            .I(N__32041));
    CEMux I__7292 (
            .O(N__32050),
            .I(N__32038));
    LocalMux I__7291 (
            .O(N__32047),
            .I(N__32035));
    Span4Mux_h I__7290 (
            .O(N__32044),
            .I(N__32032));
    Span4Mux_v I__7289 (
            .O(N__32041),
            .I(N__32029));
    LocalMux I__7288 (
            .O(N__32038),
            .I(N__32026));
    Span4Mux_h I__7287 (
            .O(N__32035),
            .I(N__32023));
    Span4Mux_v I__7286 (
            .O(N__32032),
            .I(N__32016));
    Span4Mux_h I__7285 (
            .O(N__32029),
            .I(N__32016));
    Span4Mux_v I__7284 (
            .O(N__32026),
            .I(N__32016));
    Odrv4 I__7283 (
            .O(N__32023),
            .I(\this_ppu.N_756_0_0 ));
    Odrv4 I__7282 (
            .O(N__32016),
            .I(\this_ppu.N_756_0_0 ));
    InMux I__7281 (
            .O(N__32011),
            .I(N__32008));
    LocalMux I__7280 (
            .O(N__32008),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__7279 (
            .O(N__32005),
            .I(N__32002));
    LocalMux I__7278 (
            .O(N__32002),
            .I(N__31999));
    Span4Mux_h I__7277 (
            .O(N__31999),
            .I(N__31996));
    Odrv4 I__7276 (
            .O(N__31996),
            .I(M_this_oam_ram_write_data_2));
    InMux I__7275 (
            .O(N__31993),
            .I(N__31990));
    LocalMux I__7274 (
            .O(N__31990),
            .I(N__31987));
    Span4Mux_v I__7273 (
            .O(N__31987),
            .I(N__31984));
    Span4Mux_h I__7272 (
            .O(N__31984),
            .I(N__31981));
    Odrv4 I__7271 (
            .O(N__31981),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__7270 (
            .O(N__31978),
            .I(N__31975));
    LocalMux I__7269 (
            .O(N__31975),
            .I(N__31972));
    Span4Mux_h I__7268 (
            .O(N__31972),
            .I(N__31969));
    Odrv4 I__7267 (
            .O(N__31969),
            .I(M_this_oam_ram_write_data_16));
    InMux I__7266 (
            .O(N__31966),
            .I(N__31963));
    LocalMux I__7265 (
            .O(N__31963),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__7264 (
            .O(N__31960),
            .I(N__31957));
    LocalMux I__7263 (
            .O(N__31957),
            .I(N__31954));
    Span4Mux_v I__7262 (
            .O(N__31954),
            .I(N__31951));
    Odrv4 I__7261 (
            .O(N__31951),
            .I(M_this_oam_ram_write_data_5));
    InMux I__7260 (
            .O(N__31948),
            .I(N__31945));
    LocalMux I__7259 (
            .O(N__31945),
            .I(N__31942));
    Odrv4 I__7258 (
            .O(N__31942),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__7257 (
            .O(N__31939),
            .I(N__31936));
    LocalMux I__7256 (
            .O(N__31936),
            .I(N__31933));
    Odrv12 I__7255 (
            .O(N__31933),
            .I(M_this_oam_ram_write_data_15));
    InMux I__7254 (
            .O(N__31930),
            .I(N__31927));
    LocalMux I__7253 (
            .O(N__31927),
            .I(M_this_data_tmp_qZ0Z_19));
    InMux I__7252 (
            .O(N__31924),
            .I(N__31921));
    LocalMux I__7251 (
            .O(N__31921),
            .I(N__31918));
    Span4Mux_h I__7250 (
            .O(N__31918),
            .I(N__31915));
    Odrv4 I__7249 (
            .O(N__31915),
            .I(M_this_oam_ram_write_data_19));
    CascadeMux I__7248 (
            .O(N__31912),
            .I(N__31909));
    InMux I__7247 (
            .O(N__31909),
            .I(N__31906));
    LocalMux I__7246 (
            .O(N__31906),
            .I(\this_ppu.M_oam_cache_read_data_i_17 ));
    InMux I__7245 (
            .O(N__31903),
            .I(N__31900));
    LocalMux I__7244 (
            .O(N__31900),
            .I(N__31897));
    Span4Mux_h I__7243 (
            .O(N__31897),
            .I(N__31894));
    Odrv4 I__7242 (
            .O(N__31894),
            .I(\this_ppu.oam_cache.mem_17 ));
    InMux I__7241 (
            .O(N__31891),
            .I(N__31888));
    LocalMux I__7240 (
            .O(N__31888),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_17 ));
    CascadeMux I__7239 (
            .O(N__31885),
            .I(N__31881));
    InMux I__7238 (
            .O(N__31884),
            .I(N__31877));
    InMux I__7237 (
            .O(N__31881),
            .I(N__31873));
    InMux I__7236 (
            .O(N__31880),
            .I(N__31870));
    LocalMux I__7235 (
            .O(N__31877),
            .I(N__31867));
    InMux I__7234 (
            .O(N__31876),
            .I(N__31864));
    LocalMux I__7233 (
            .O(N__31873),
            .I(N__31853));
    LocalMux I__7232 (
            .O(N__31870),
            .I(N__31853));
    Span4Mux_h I__7231 (
            .O(N__31867),
            .I(N__31853));
    LocalMux I__7230 (
            .O(N__31864),
            .I(N__31853));
    CascadeMux I__7229 (
            .O(N__31863),
            .I(N__31850));
    InMux I__7228 (
            .O(N__31862),
            .I(N__31847));
    Span4Mux_v I__7227 (
            .O(N__31853),
            .I(N__31844));
    InMux I__7226 (
            .O(N__31850),
            .I(N__31840));
    LocalMux I__7225 (
            .O(N__31847),
            .I(N__31837));
    Span4Mux_h I__7224 (
            .O(N__31844),
            .I(N__31834));
    CascadeMux I__7223 (
            .O(N__31843),
            .I(N__31831));
    LocalMux I__7222 (
            .O(N__31840),
            .I(N__31828));
    Span4Mux_v I__7221 (
            .O(N__31837),
            .I(N__31823));
    Span4Mux_h I__7220 (
            .O(N__31834),
            .I(N__31823));
    InMux I__7219 (
            .O(N__31831),
            .I(N__31820));
    Span12Mux_s11_h I__7218 (
            .O(N__31828),
            .I(N__31817));
    Span4Mux_v I__7217 (
            .O(N__31823),
            .I(N__31814));
    LocalMux I__7216 (
            .O(N__31820),
            .I(M_this_ppu_vram_addr_7));
    Odrv12 I__7215 (
            .O(N__31817),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__7214 (
            .O(N__31814),
            .I(M_this_ppu_vram_addr_7));
    InMux I__7213 (
            .O(N__31807),
            .I(N__31803));
    InMux I__7212 (
            .O(N__31806),
            .I(N__31800));
    LocalMux I__7211 (
            .O(N__31803),
            .I(N__31794));
    LocalMux I__7210 (
            .O(N__31800),
            .I(N__31794));
    InMux I__7209 (
            .O(N__31799),
            .I(N__31791));
    Span4Mux_v I__7208 (
            .O(N__31794),
            .I(N__31787));
    LocalMux I__7207 (
            .O(N__31791),
            .I(N__31784));
    InMux I__7206 (
            .O(N__31790),
            .I(N__31781));
    Sp12to4 I__7205 (
            .O(N__31787),
            .I(N__31776));
    Span12Mux_s10_v I__7204 (
            .O(N__31784),
            .I(N__31776));
    LocalMux I__7203 (
            .O(N__31781),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    Odrv12 I__7202 (
            .O(N__31776),
            .I(\this_ppu.M_vaddress_qZ0Z_1 ));
    InMux I__7201 (
            .O(N__31771),
            .I(\this_ppu.un1_M_voffset_d_cry_0 ));
    InMux I__7200 (
            .O(N__31768),
            .I(N__31759));
    InMux I__7199 (
            .O(N__31767),
            .I(N__31759));
    InMux I__7198 (
            .O(N__31766),
            .I(N__31759));
    LocalMux I__7197 (
            .O(N__31759),
            .I(N__31754));
    InMux I__7196 (
            .O(N__31758),
            .I(N__31751));
    InMux I__7195 (
            .O(N__31757),
            .I(N__31748));
    Odrv4 I__7194 (
            .O(N__31754),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7193 (
            .O(N__31751),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    LocalMux I__7192 (
            .O(N__31748),
            .I(\this_ppu.M_vaddress_qZ0Z_2 ));
    InMux I__7191 (
            .O(N__31741),
            .I(\this_ppu.un1_M_voffset_d_cry_1 ));
    CascadeMux I__7190 (
            .O(N__31738),
            .I(N__31735));
    InMux I__7189 (
            .O(N__31735),
            .I(N__31731));
    InMux I__7188 (
            .O(N__31734),
            .I(N__31728));
    LocalMux I__7187 (
            .O(N__31731),
            .I(N__31722));
    LocalMux I__7186 (
            .O(N__31728),
            .I(N__31722));
    CascadeMux I__7185 (
            .O(N__31727),
            .I(N__31719));
    Span12Mux_s10_v I__7184 (
            .O(N__31722),
            .I(N__31713));
    InMux I__7183 (
            .O(N__31719),
            .I(N__31708));
    InMux I__7182 (
            .O(N__31718),
            .I(N__31708));
    InMux I__7181 (
            .O(N__31717),
            .I(N__31705));
    InMux I__7180 (
            .O(N__31716),
            .I(N__31702));
    Span12Mux_v I__7179 (
            .O(N__31713),
            .I(N__31699));
    LocalMux I__7178 (
            .O(N__31708),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    LocalMux I__7177 (
            .O(N__31705),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    LocalMux I__7176 (
            .O(N__31702),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    Odrv12 I__7175 (
            .O(N__31699),
            .I(\this_ppu.M_vaddress_qZ0Z_3 ));
    InMux I__7174 (
            .O(N__31690),
            .I(\this_ppu.un1_M_voffset_d_cry_2 ));
    CascadeMux I__7173 (
            .O(N__31687),
            .I(N__31684));
    InMux I__7172 (
            .O(N__31684),
            .I(N__31681));
    LocalMux I__7171 (
            .O(N__31681),
            .I(N__31678));
    Span4Mux_h I__7170 (
            .O(N__31678),
            .I(N__31674));
    CascadeMux I__7169 (
            .O(N__31677),
            .I(N__31670));
    Sp12to4 I__7168 (
            .O(N__31674),
            .I(N__31666));
    InMux I__7167 (
            .O(N__31673),
            .I(N__31663));
    InMux I__7166 (
            .O(N__31670),
            .I(N__31660));
    InMux I__7165 (
            .O(N__31669),
            .I(N__31657));
    Span12Mux_v I__7164 (
            .O(N__31666),
            .I(N__31654));
    LocalMux I__7163 (
            .O(N__31663),
            .I(\this_ppu.M_vaddress_qZ0Z_4 ));
    LocalMux I__7162 (
            .O(N__31660),
            .I(\this_ppu.M_vaddress_qZ0Z_4 ));
    LocalMux I__7161 (
            .O(N__31657),
            .I(\this_ppu.M_vaddress_qZ0Z_4 ));
    Odrv12 I__7160 (
            .O(N__31654),
            .I(\this_ppu.M_vaddress_qZ0Z_4 ));
    InMux I__7159 (
            .O(N__31645),
            .I(\this_ppu.un1_M_voffset_d_cry_3 ));
    CascadeMux I__7158 (
            .O(N__31642),
            .I(N__31639));
    InMux I__7157 (
            .O(N__31639),
            .I(N__31636));
    LocalMux I__7156 (
            .O(N__31636),
            .I(N__31633));
    Span4Mux_h I__7155 (
            .O(N__31633),
            .I(N__31628));
    CascadeMux I__7154 (
            .O(N__31632),
            .I(N__31625));
    CascadeMux I__7153 (
            .O(N__31631),
            .I(N__31622));
    Sp12to4 I__7152 (
            .O(N__31628),
            .I(N__31618));
    InMux I__7151 (
            .O(N__31625),
            .I(N__31610));
    InMux I__7150 (
            .O(N__31622),
            .I(N__31610));
    InMux I__7149 (
            .O(N__31621),
            .I(N__31610));
    Span12Mux_v I__7148 (
            .O(N__31618),
            .I(N__31607));
    InMux I__7147 (
            .O(N__31617),
            .I(N__31604));
    LocalMux I__7146 (
            .O(N__31610),
            .I(\this_ppu.M_vaddress_qZ0Z_5 ));
    Odrv12 I__7145 (
            .O(N__31607),
            .I(\this_ppu.M_vaddress_qZ0Z_5 ));
    LocalMux I__7144 (
            .O(N__31604),
            .I(\this_ppu.M_vaddress_qZ0Z_5 ));
    InMux I__7143 (
            .O(N__31597),
            .I(\this_ppu.un1_M_voffset_d_cry_4 ));
    CascadeMux I__7142 (
            .O(N__31594),
            .I(N__31591));
    InMux I__7141 (
            .O(N__31591),
            .I(N__31588));
    LocalMux I__7140 (
            .O(N__31588),
            .I(N__31585));
    Span4Mux_v I__7139 (
            .O(N__31585),
            .I(N__31582));
    Span4Mux_h I__7138 (
            .O(N__31582),
            .I(N__31578));
    CascadeMux I__7137 (
            .O(N__31581),
            .I(N__31573));
    Sp12to4 I__7136 (
            .O(N__31578),
            .I(N__31570));
    InMux I__7135 (
            .O(N__31577),
            .I(N__31565));
    InMux I__7134 (
            .O(N__31576),
            .I(N__31565));
    InMux I__7133 (
            .O(N__31573),
            .I(N__31562));
    Span12Mux_v I__7132 (
            .O(N__31570),
            .I(N__31559));
    LocalMux I__7131 (
            .O(N__31565),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    LocalMux I__7130 (
            .O(N__31562),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    Odrv12 I__7129 (
            .O(N__31559),
            .I(\this_ppu.M_vaddress_qZ0Z_6 ));
    InMux I__7128 (
            .O(N__31552),
            .I(\this_ppu.un1_oam_data_1_cry_8 ));
    InMux I__7127 (
            .O(N__31549),
            .I(N__31545));
    InMux I__7126 (
            .O(N__31548),
            .I(N__31542));
    LocalMux I__7125 (
            .O(N__31545),
            .I(N__31539));
    LocalMux I__7124 (
            .O(N__31542),
            .I(N__31535));
    Span4Mux_v I__7123 (
            .O(N__31539),
            .I(N__31532));
    InMux I__7122 (
            .O(N__31538),
            .I(N__31529));
    Odrv4 I__7121 (
            .O(N__31535),
            .I(\this_ppu.un1_oam_data_1_cry_8_THRU_CO ));
    Odrv4 I__7120 (
            .O(N__31532),
            .I(\this_ppu.un1_oam_data_1_cry_8_THRU_CO ));
    LocalMux I__7119 (
            .O(N__31529),
            .I(\this_ppu.un1_oam_data_1_cry_8_THRU_CO ));
    CascadeMux I__7118 (
            .O(N__31522),
            .I(N__31519));
    InMux I__7117 (
            .O(N__31519),
            .I(N__31516));
    LocalMux I__7116 (
            .O(N__31516),
            .I(\this_ppu.vspr_cry_0_c_inv_RNIFK43 ));
    CascadeMux I__7115 (
            .O(N__31513),
            .I(N__31509));
    CascadeMux I__7114 (
            .O(N__31512),
            .I(N__31506));
    InMux I__7113 (
            .O(N__31509),
            .I(N__31500));
    InMux I__7112 (
            .O(N__31506),
            .I(N__31497));
    CascadeMux I__7111 (
            .O(N__31505),
            .I(N__31494));
    CascadeMux I__7110 (
            .O(N__31504),
            .I(N__31490));
    CascadeMux I__7109 (
            .O(N__31503),
            .I(N__31487));
    LocalMux I__7108 (
            .O(N__31500),
            .I(N__31480));
    LocalMux I__7107 (
            .O(N__31497),
            .I(N__31480));
    InMux I__7106 (
            .O(N__31494),
            .I(N__31477));
    CascadeMux I__7105 (
            .O(N__31493),
            .I(N__31474));
    InMux I__7104 (
            .O(N__31490),
            .I(N__31470));
    InMux I__7103 (
            .O(N__31487),
            .I(N__31467));
    CascadeMux I__7102 (
            .O(N__31486),
            .I(N__31464));
    CascadeMux I__7101 (
            .O(N__31485),
            .I(N__31461));
    Span4Mux_s2_v I__7100 (
            .O(N__31480),
            .I(N__31454));
    LocalMux I__7099 (
            .O(N__31477),
            .I(N__31454));
    InMux I__7098 (
            .O(N__31474),
            .I(N__31451));
    CascadeMux I__7097 (
            .O(N__31473),
            .I(N__31448));
    LocalMux I__7096 (
            .O(N__31470),
            .I(N__31442));
    LocalMux I__7095 (
            .O(N__31467),
            .I(N__31442));
    InMux I__7094 (
            .O(N__31464),
            .I(N__31439));
    InMux I__7093 (
            .O(N__31461),
            .I(N__31436));
    CascadeMux I__7092 (
            .O(N__31460),
            .I(N__31433));
    CascadeMux I__7091 (
            .O(N__31459),
            .I(N__31430));
    Span4Mux_v I__7090 (
            .O(N__31454),
            .I(N__31424));
    LocalMux I__7089 (
            .O(N__31451),
            .I(N__31424));
    InMux I__7088 (
            .O(N__31448),
            .I(N__31421));
    CascadeMux I__7087 (
            .O(N__31447),
            .I(N__31418));
    Span4Mux_v I__7086 (
            .O(N__31442),
            .I(N__31410));
    LocalMux I__7085 (
            .O(N__31439),
            .I(N__31410));
    LocalMux I__7084 (
            .O(N__31436),
            .I(N__31410));
    InMux I__7083 (
            .O(N__31433),
            .I(N__31407));
    InMux I__7082 (
            .O(N__31430),
            .I(N__31404));
    CascadeMux I__7081 (
            .O(N__31429),
            .I(N__31401));
    Span4Mux_v I__7080 (
            .O(N__31424),
            .I(N__31395));
    LocalMux I__7079 (
            .O(N__31421),
            .I(N__31395));
    InMux I__7078 (
            .O(N__31418),
            .I(N__31392));
    CascadeMux I__7077 (
            .O(N__31417),
            .I(N__31389));
    Span4Mux_v I__7076 (
            .O(N__31410),
            .I(N__31381));
    LocalMux I__7075 (
            .O(N__31407),
            .I(N__31381));
    LocalMux I__7074 (
            .O(N__31404),
            .I(N__31381));
    InMux I__7073 (
            .O(N__31401),
            .I(N__31378));
    CascadeMux I__7072 (
            .O(N__31400),
            .I(N__31375));
    Span4Mux_v I__7071 (
            .O(N__31395),
            .I(N__31370));
    LocalMux I__7070 (
            .O(N__31392),
            .I(N__31370));
    InMux I__7069 (
            .O(N__31389),
            .I(N__31367));
    CascadeMux I__7068 (
            .O(N__31388),
            .I(N__31364));
    Sp12to4 I__7067 (
            .O(N__31381),
            .I(N__31361));
    LocalMux I__7066 (
            .O(N__31378),
            .I(N__31358));
    InMux I__7065 (
            .O(N__31375),
            .I(N__31355));
    Span4Mux_h I__7064 (
            .O(N__31370),
            .I(N__31350));
    LocalMux I__7063 (
            .O(N__31367),
            .I(N__31350));
    InMux I__7062 (
            .O(N__31364),
            .I(N__31347));
    Span12Mux_v I__7061 (
            .O(N__31361),
            .I(N__31344));
    Span12Mux_s11_h I__7060 (
            .O(N__31358),
            .I(N__31341));
    LocalMux I__7059 (
            .O(N__31355),
            .I(N__31338));
    Span4Mux_v I__7058 (
            .O(N__31350),
            .I(N__31333));
    LocalMux I__7057 (
            .O(N__31347),
            .I(N__31333));
    Span12Mux_h I__7056 (
            .O(N__31344),
            .I(N__31328));
    Span12Mux_v I__7055 (
            .O(N__31341),
            .I(N__31328));
    Span12Mux_s11_h I__7054 (
            .O(N__31338),
            .I(N__31325));
    Span4Mux_h I__7053 (
            .O(N__31333),
            .I(N__31322));
    Odrv12 I__7052 (
            .O(N__31328),
            .I(M_this_ppu_spr_addr_4));
    Odrv12 I__7051 (
            .O(N__31325),
            .I(M_this_ppu_spr_addr_4));
    Odrv4 I__7050 (
            .O(N__31322),
            .I(M_this_ppu_spr_addr_4));
    InMux I__7049 (
            .O(N__31315),
            .I(\this_ppu.vspr_cry_0 ));
    InMux I__7048 (
            .O(N__31312),
            .I(\this_ppu.vspr_cry_1 ));
    CascadeMux I__7047 (
            .O(N__31309),
            .I(N__31305));
    CascadeMux I__7046 (
            .O(N__31308),
            .I(N__31302));
    InMux I__7045 (
            .O(N__31305),
            .I(N__31298));
    InMux I__7044 (
            .O(N__31302),
            .I(N__31295));
    CascadeMux I__7043 (
            .O(N__31301),
            .I(N__31292));
    LocalMux I__7042 (
            .O(N__31298),
            .I(N__31286));
    LocalMux I__7041 (
            .O(N__31295),
            .I(N__31286));
    InMux I__7040 (
            .O(N__31292),
            .I(N__31283));
    CascadeMux I__7039 (
            .O(N__31291),
            .I(N__31280));
    Span4Mux_s2_v I__7038 (
            .O(N__31286),
            .I(N__31272));
    LocalMux I__7037 (
            .O(N__31283),
            .I(N__31272));
    InMux I__7036 (
            .O(N__31280),
            .I(N__31269));
    CascadeMux I__7035 (
            .O(N__31279),
            .I(N__31266));
    CascadeMux I__7034 (
            .O(N__31278),
            .I(N__31262));
    CascadeMux I__7033 (
            .O(N__31277),
            .I(N__31259));
    Span4Mux_v I__7032 (
            .O(N__31272),
            .I(N__31252));
    LocalMux I__7031 (
            .O(N__31269),
            .I(N__31252));
    InMux I__7030 (
            .O(N__31266),
            .I(N__31249));
    CascadeMux I__7029 (
            .O(N__31265),
            .I(N__31246));
    InMux I__7028 (
            .O(N__31262),
            .I(N__31242));
    InMux I__7027 (
            .O(N__31259),
            .I(N__31239));
    CascadeMux I__7026 (
            .O(N__31258),
            .I(N__31236));
    CascadeMux I__7025 (
            .O(N__31257),
            .I(N__31233));
    Span4Mux_h I__7024 (
            .O(N__31252),
            .I(N__31226));
    LocalMux I__7023 (
            .O(N__31249),
            .I(N__31226));
    InMux I__7022 (
            .O(N__31246),
            .I(N__31223));
    CascadeMux I__7021 (
            .O(N__31245),
            .I(N__31220));
    LocalMux I__7020 (
            .O(N__31242),
            .I(N__31214));
    LocalMux I__7019 (
            .O(N__31239),
            .I(N__31214));
    InMux I__7018 (
            .O(N__31236),
            .I(N__31211));
    InMux I__7017 (
            .O(N__31233),
            .I(N__31208));
    CascadeMux I__7016 (
            .O(N__31232),
            .I(N__31205));
    CascadeMux I__7015 (
            .O(N__31231),
            .I(N__31202));
    Span4Mux_v I__7014 (
            .O(N__31226),
            .I(N__31197));
    LocalMux I__7013 (
            .O(N__31223),
            .I(N__31197));
    InMux I__7012 (
            .O(N__31220),
            .I(N__31194));
    CascadeMux I__7011 (
            .O(N__31219),
            .I(N__31191));
    Span4Mux_v I__7010 (
            .O(N__31214),
            .I(N__31183));
    LocalMux I__7009 (
            .O(N__31211),
            .I(N__31183));
    LocalMux I__7008 (
            .O(N__31208),
            .I(N__31183));
    InMux I__7007 (
            .O(N__31205),
            .I(N__31180));
    InMux I__7006 (
            .O(N__31202),
            .I(N__31177));
    Span4Mux_h I__7005 (
            .O(N__31197),
            .I(N__31172));
    LocalMux I__7004 (
            .O(N__31194),
            .I(N__31172));
    InMux I__7003 (
            .O(N__31191),
            .I(N__31169));
    CascadeMux I__7002 (
            .O(N__31190),
            .I(N__31166));
    Span4Mux_v I__7001 (
            .O(N__31183),
            .I(N__31158));
    LocalMux I__7000 (
            .O(N__31180),
            .I(N__31158));
    LocalMux I__6999 (
            .O(N__31177),
            .I(N__31158));
    Span4Mux_v I__6998 (
            .O(N__31172),
            .I(N__31153));
    LocalMux I__6997 (
            .O(N__31169),
            .I(N__31153));
    InMux I__6996 (
            .O(N__31166),
            .I(N__31150));
    CascadeMux I__6995 (
            .O(N__31165),
            .I(N__31147));
    Sp12to4 I__6994 (
            .O(N__31158),
            .I(N__31144));
    Span4Mux_h I__6993 (
            .O(N__31153),
            .I(N__31139));
    LocalMux I__6992 (
            .O(N__31150),
            .I(N__31139));
    InMux I__6991 (
            .O(N__31147),
            .I(N__31136));
    Span12Mux_v I__6990 (
            .O(N__31144),
            .I(N__31133));
    Span4Mux_v I__6989 (
            .O(N__31139),
            .I(N__31128));
    LocalMux I__6988 (
            .O(N__31136),
            .I(N__31128));
    Span12Mux_h I__6987 (
            .O(N__31133),
            .I(N__31125));
    Span4Mux_h I__6986 (
            .O(N__31128),
            .I(N__31122));
    Odrv12 I__6985 (
            .O(N__31125),
            .I(M_this_ppu_spr_addr_5));
    Odrv4 I__6984 (
            .O(N__31122),
            .I(M_this_ppu_spr_addr_5));
    InMux I__6983 (
            .O(N__31117),
            .I(N__31114));
    LocalMux I__6982 (
            .O(N__31114),
            .I(\this_ppu.M_hoffset_q_i_8 ));
    InMux I__6981 (
            .O(N__31111),
            .I(\this_ppu.un1_M_hoffset_q_2_cry_8 ));
    InMux I__6980 (
            .O(N__31108),
            .I(N__31105));
    LocalMux I__6979 (
            .O(N__31105),
            .I(\this_ppu.vspr12_0 ));
    InMux I__6978 (
            .O(N__31102),
            .I(N__31099));
    LocalMux I__6977 (
            .O(N__31099),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0 ));
    CascadeMux I__6976 (
            .O(N__31096),
            .I(N__31092));
    CascadeMux I__6975 (
            .O(N__31095),
            .I(N__31089));
    InMux I__6974 (
            .O(N__31092),
            .I(N__31083));
    InMux I__6973 (
            .O(N__31089),
            .I(N__31080));
    CascadeMux I__6972 (
            .O(N__31088),
            .I(N__31077));
    CascadeMux I__6971 (
            .O(N__31087),
            .I(N__31073));
    CascadeMux I__6970 (
            .O(N__31086),
            .I(N__31070));
    LocalMux I__6969 (
            .O(N__31083),
            .I(N__31064));
    LocalMux I__6968 (
            .O(N__31080),
            .I(N__31064));
    InMux I__6967 (
            .O(N__31077),
            .I(N__31061));
    CascadeMux I__6966 (
            .O(N__31076),
            .I(N__31058));
    InMux I__6965 (
            .O(N__31073),
            .I(N__31054));
    InMux I__6964 (
            .O(N__31070),
            .I(N__31051));
    CascadeMux I__6963 (
            .O(N__31069),
            .I(N__31048));
    Span4Mux_s2_v I__6962 (
            .O(N__31064),
            .I(N__31042));
    LocalMux I__6961 (
            .O(N__31061),
            .I(N__31042));
    InMux I__6960 (
            .O(N__31058),
            .I(N__31039));
    CascadeMux I__6959 (
            .O(N__31057),
            .I(N__31036));
    LocalMux I__6958 (
            .O(N__31054),
            .I(N__31032));
    LocalMux I__6957 (
            .O(N__31051),
            .I(N__31029));
    InMux I__6956 (
            .O(N__31048),
            .I(N__31026));
    CascadeMux I__6955 (
            .O(N__31047),
            .I(N__31023));
    Span4Mux_v I__6954 (
            .O(N__31042),
            .I(N__31017));
    LocalMux I__6953 (
            .O(N__31039),
            .I(N__31017));
    InMux I__6952 (
            .O(N__31036),
            .I(N__31014));
    CascadeMux I__6951 (
            .O(N__31035),
            .I(N__31011));
    Span4Mux_v I__6950 (
            .O(N__31032),
            .I(N__31002));
    Span4Mux_h I__6949 (
            .O(N__31029),
            .I(N__31002));
    LocalMux I__6948 (
            .O(N__31026),
            .I(N__31002));
    InMux I__6947 (
            .O(N__31023),
            .I(N__30999));
    CascadeMux I__6946 (
            .O(N__31022),
            .I(N__30996));
    Span4Mux_h I__6945 (
            .O(N__31017),
            .I(N__30990));
    LocalMux I__6944 (
            .O(N__31014),
            .I(N__30990));
    InMux I__6943 (
            .O(N__31011),
            .I(N__30987));
    CascadeMux I__6942 (
            .O(N__31010),
            .I(N__30984));
    CascadeMux I__6941 (
            .O(N__31009),
            .I(N__30980));
    Span4Mux_v I__6940 (
            .O(N__31002),
            .I(N__30975));
    LocalMux I__6939 (
            .O(N__30999),
            .I(N__30975));
    InMux I__6938 (
            .O(N__30996),
            .I(N__30972));
    CascadeMux I__6937 (
            .O(N__30995),
            .I(N__30969));
    Span4Mux_v I__6936 (
            .O(N__30990),
            .I(N__30964));
    LocalMux I__6935 (
            .O(N__30987),
            .I(N__30964));
    InMux I__6934 (
            .O(N__30984),
            .I(N__30961));
    CascadeMux I__6933 (
            .O(N__30983),
            .I(N__30958));
    InMux I__6932 (
            .O(N__30980),
            .I(N__30955));
    Span4Mux_h I__6931 (
            .O(N__30975),
            .I(N__30950));
    LocalMux I__6930 (
            .O(N__30972),
            .I(N__30950));
    InMux I__6929 (
            .O(N__30969),
            .I(N__30946));
    Span4Mux_h I__6928 (
            .O(N__30964),
            .I(N__30941));
    LocalMux I__6927 (
            .O(N__30961),
            .I(N__30941));
    InMux I__6926 (
            .O(N__30958),
            .I(N__30938));
    LocalMux I__6925 (
            .O(N__30955),
            .I(N__30935));
    Span4Mux_v I__6924 (
            .O(N__30950),
            .I(N__30932));
    CascadeMux I__6923 (
            .O(N__30949),
            .I(N__30929));
    LocalMux I__6922 (
            .O(N__30946),
            .I(N__30926));
    Span4Mux_v I__6921 (
            .O(N__30941),
            .I(N__30921));
    LocalMux I__6920 (
            .O(N__30938),
            .I(N__30921));
    Span12Mux_h I__6919 (
            .O(N__30935),
            .I(N__30918));
    Sp12to4 I__6918 (
            .O(N__30932),
            .I(N__30915));
    InMux I__6917 (
            .O(N__30929),
            .I(N__30912));
    Span4Mux_h I__6916 (
            .O(N__30926),
            .I(N__30907));
    Span4Mux_h I__6915 (
            .O(N__30921),
            .I(N__30907));
    Span12Mux_v I__6914 (
            .O(N__30918),
            .I(N__30900));
    Span12Mux_h I__6913 (
            .O(N__30915),
            .I(N__30900));
    LocalMux I__6912 (
            .O(N__30912),
            .I(N__30900));
    Odrv4 I__6911 (
            .O(N__30907),
            .I(M_this_ppu_spr_addr_1));
    Odrv12 I__6910 (
            .O(N__30900),
            .I(M_this_ppu_spr_addr_1));
    InMux I__6909 (
            .O(N__30895),
            .I(\this_ppu.hspr_cry_0 ));
    InMux I__6908 (
            .O(N__30892),
            .I(\this_ppu.hspr_cry_1 ));
    CascadeMux I__6907 (
            .O(N__30889),
            .I(N__30885));
    CascadeMux I__6906 (
            .O(N__30888),
            .I(N__30882));
    InMux I__6905 (
            .O(N__30885),
            .I(N__30876));
    InMux I__6904 (
            .O(N__30882),
            .I(N__30873));
    CascadeMux I__6903 (
            .O(N__30881),
            .I(N__30870));
    CascadeMux I__6902 (
            .O(N__30880),
            .I(N__30867));
    CascadeMux I__6901 (
            .O(N__30879),
            .I(N__30863));
    LocalMux I__6900 (
            .O(N__30876),
            .I(N__30859));
    LocalMux I__6899 (
            .O(N__30873),
            .I(N__30856));
    InMux I__6898 (
            .O(N__30870),
            .I(N__30853));
    InMux I__6897 (
            .O(N__30867),
            .I(N__30850));
    CascadeMux I__6896 (
            .O(N__30866),
            .I(N__30847));
    InMux I__6895 (
            .O(N__30863),
            .I(N__30844));
    CascadeMux I__6894 (
            .O(N__30862),
            .I(N__30841));
    Span4Mux_v I__6893 (
            .O(N__30859),
            .I(N__30832));
    Span4Mux_h I__6892 (
            .O(N__30856),
            .I(N__30832));
    LocalMux I__6891 (
            .O(N__30853),
            .I(N__30832));
    LocalMux I__6890 (
            .O(N__30850),
            .I(N__30829));
    InMux I__6889 (
            .O(N__30847),
            .I(N__30826));
    LocalMux I__6888 (
            .O(N__30844),
            .I(N__30823));
    InMux I__6887 (
            .O(N__30841),
            .I(N__30820));
    CascadeMux I__6886 (
            .O(N__30840),
            .I(N__30817));
    CascadeMux I__6885 (
            .O(N__30839),
            .I(N__30812));
    Span4Mux_v I__6884 (
            .O(N__30832),
            .I(N__30803));
    Span4Mux_h I__6883 (
            .O(N__30829),
            .I(N__30803));
    LocalMux I__6882 (
            .O(N__30826),
            .I(N__30803));
    Span4Mux_s0_v I__6881 (
            .O(N__30823),
            .I(N__30797));
    LocalMux I__6880 (
            .O(N__30820),
            .I(N__30797));
    InMux I__6879 (
            .O(N__30817),
            .I(N__30794));
    CascadeMux I__6878 (
            .O(N__30816),
            .I(N__30791));
    CascadeMux I__6877 (
            .O(N__30815),
            .I(N__30788));
    InMux I__6876 (
            .O(N__30812),
            .I(N__30784));
    CascadeMux I__6875 (
            .O(N__30811),
            .I(N__30781));
    CascadeMux I__6874 (
            .O(N__30810),
            .I(N__30778));
    Span4Mux_v I__6873 (
            .O(N__30803),
            .I(N__30775));
    CascadeMux I__6872 (
            .O(N__30802),
            .I(N__30772));
    Span4Mux_v I__6871 (
            .O(N__30797),
            .I(N__30769));
    LocalMux I__6870 (
            .O(N__30794),
            .I(N__30766));
    InMux I__6869 (
            .O(N__30791),
            .I(N__30763));
    InMux I__6868 (
            .O(N__30788),
            .I(N__30760));
    CascadeMux I__6867 (
            .O(N__30787),
            .I(N__30757));
    LocalMux I__6866 (
            .O(N__30784),
            .I(N__30754));
    InMux I__6865 (
            .O(N__30781),
            .I(N__30751));
    InMux I__6864 (
            .O(N__30778),
            .I(N__30747));
    Span4Mux_h I__6863 (
            .O(N__30775),
            .I(N__30744));
    InMux I__6862 (
            .O(N__30772),
            .I(N__30741));
    Span4Mux_v I__6861 (
            .O(N__30769),
            .I(N__30734));
    Span4Mux_h I__6860 (
            .O(N__30766),
            .I(N__30734));
    LocalMux I__6859 (
            .O(N__30763),
            .I(N__30734));
    LocalMux I__6858 (
            .O(N__30760),
            .I(N__30731));
    InMux I__6857 (
            .O(N__30757),
            .I(N__30728));
    Span12Mux_h I__6856 (
            .O(N__30754),
            .I(N__30723));
    LocalMux I__6855 (
            .O(N__30751),
            .I(N__30723));
    CascadeMux I__6854 (
            .O(N__30750),
            .I(N__30720));
    LocalMux I__6853 (
            .O(N__30747),
            .I(N__30717));
    Span4Mux_h I__6852 (
            .O(N__30744),
            .I(N__30714));
    LocalMux I__6851 (
            .O(N__30741),
            .I(N__30711));
    Span4Mux_v I__6850 (
            .O(N__30734),
            .I(N__30704));
    Span4Mux_h I__6849 (
            .O(N__30731),
            .I(N__30704));
    LocalMux I__6848 (
            .O(N__30728),
            .I(N__30704));
    Span12Mux_h I__6847 (
            .O(N__30723),
            .I(N__30701));
    InMux I__6846 (
            .O(N__30720),
            .I(N__30698));
    Span12Mux_s11_h I__6845 (
            .O(N__30717),
            .I(N__30695));
    Span4Mux_h I__6844 (
            .O(N__30714),
            .I(N__30688));
    Span4Mux_v I__6843 (
            .O(N__30711),
            .I(N__30688));
    Span4Mux_v I__6842 (
            .O(N__30704),
            .I(N__30688));
    Span12Mux_v I__6841 (
            .O(N__30701),
            .I(N__30683));
    LocalMux I__6840 (
            .O(N__30698),
            .I(N__30683));
    Odrv12 I__6839 (
            .O(N__30695),
            .I(M_this_ppu_spr_addr_2));
    Odrv4 I__6838 (
            .O(N__30688),
            .I(M_this_ppu_spr_addr_2));
    Odrv12 I__6837 (
            .O(N__30683),
            .I(M_this_ppu_spr_addr_2));
    CascadeMux I__6836 (
            .O(N__30676),
            .I(N__30673));
    InMux I__6835 (
            .O(N__30673),
            .I(N__30670));
    LocalMux I__6834 (
            .O(N__30670),
            .I(\this_ppu.M_oam_cache_read_data_i_9 ));
    CascadeMux I__6833 (
            .O(N__30667),
            .I(\this_ppu.N_424_cascade_ ));
    InMux I__6832 (
            .O(N__30664),
            .I(N__30661));
    LocalMux I__6831 (
            .O(N__30661),
            .I(N__30658));
    Odrv4 I__6830 (
            .O(N__30658),
            .I(\this_ppu.N_449 ));
    InMux I__6829 (
            .O(N__30655),
            .I(N__30652));
    LocalMux I__6828 (
            .O(N__30652),
            .I(M_this_state_q_RNI1G0LZ0Z_1));
    CascadeMux I__6827 (
            .O(N__30649),
            .I(N__30646));
    InMux I__6826 (
            .O(N__30646),
            .I(N__30640));
    InMux I__6825 (
            .O(N__30645),
            .I(N__30640));
    LocalMux I__6824 (
            .O(N__30640),
            .I(N__30637));
    Odrv4 I__6823 (
            .O(N__30637),
            .I(\this_ppu.N_341_0 ));
    InMux I__6822 (
            .O(N__30634),
            .I(N__30629));
    InMux I__6821 (
            .O(N__30633),
            .I(N__30622));
    InMux I__6820 (
            .O(N__30632),
            .I(N__30619));
    LocalMux I__6819 (
            .O(N__30629),
            .I(N__30616));
    InMux I__6818 (
            .O(N__30628),
            .I(N__30611));
    InMux I__6817 (
            .O(N__30627),
            .I(N__30611));
    InMux I__6816 (
            .O(N__30626),
            .I(N__30608));
    InMux I__6815 (
            .O(N__30625),
            .I(N__30605));
    LocalMux I__6814 (
            .O(N__30622),
            .I(N__30594));
    LocalMux I__6813 (
            .O(N__30619),
            .I(N__30594));
    Span4Mux_h I__6812 (
            .O(N__30616),
            .I(N__30594));
    LocalMux I__6811 (
            .O(N__30611),
            .I(N__30594));
    LocalMux I__6810 (
            .O(N__30608),
            .I(N__30594));
    LocalMux I__6809 (
            .O(N__30605),
            .I(N__30591));
    Span4Mux_v I__6808 (
            .O(N__30594),
            .I(N__30588));
    Span4Mux_h I__6807 (
            .O(N__30591),
            .I(N__30585));
    Span4Mux_h I__6806 (
            .O(N__30588),
            .I(N__30582));
    Odrv4 I__6805 (
            .O(N__30585),
            .I(\this_ppu.N_934 ));
    Odrv4 I__6804 (
            .O(N__30582),
            .I(\this_ppu.N_934 ));
    InMux I__6803 (
            .O(N__30577),
            .I(N__30573));
    InMux I__6802 (
            .O(N__30576),
            .I(N__30567));
    LocalMux I__6801 (
            .O(N__30573),
            .I(N__30564));
    InMux I__6800 (
            .O(N__30572),
            .I(N__30561));
    InMux I__6799 (
            .O(N__30571),
            .I(N__30556));
    InMux I__6798 (
            .O(N__30570),
            .I(N__30556));
    LocalMux I__6797 (
            .O(N__30567),
            .I(M_this_state_qZ0Z_5));
    Odrv12 I__6796 (
            .O(N__30564),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__6795 (
            .O(N__30561),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__6794 (
            .O(N__30556),
            .I(M_this_state_qZ0Z_5));
    InMux I__6793 (
            .O(N__30547),
            .I(N__30544));
    LocalMux I__6792 (
            .O(N__30544),
            .I(N__30540));
    InMux I__6791 (
            .O(N__30543),
            .I(N__30535));
    Span4Mux_h I__6790 (
            .O(N__30540),
            .I(N__30532));
    InMux I__6789 (
            .O(N__30539),
            .I(N__30529));
    InMux I__6788 (
            .O(N__30538),
            .I(N__30526));
    LocalMux I__6787 (
            .O(N__30535),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__6786 (
            .O(N__30532),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__6785 (
            .O(N__30529),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__6784 (
            .O(N__30526),
            .I(M_this_state_qZ0Z_4));
    InMux I__6783 (
            .O(N__30517),
            .I(N__30514));
    LocalMux I__6782 (
            .O(N__30514),
            .I(this_ppu_un20_i_a4_0_a2_0_a2_0_2));
    CascadeMux I__6781 (
            .O(N__30511),
            .I(N_311_0_cascade_));
    InMux I__6780 (
            .O(N__30508),
            .I(N__30505));
    LocalMux I__6779 (
            .O(N__30505),
            .I(M_this_state_q_RNI244K2Z0Z_10));
    InMux I__6778 (
            .O(N__30502),
            .I(N__30495));
    InMux I__6777 (
            .O(N__30501),
            .I(N__30491));
    InMux I__6776 (
            .O(N__30500),
            .I(N__30486));
    InMux I__6775 (
            .O(N__30499),
            .I(N__30486));
    InMux I__6774 (
            .O(N__30498),
            .I(N__30483));
    LocalMux I__6773 (
            .O(N__30495),
            .I(N__30480));
    InMux I__6772 (
            .O(N__30494),
            .I(N__30477));
    LocalMux I__6771 (
            .O(N__30491),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__6770 (
            .O(N__30486),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__6769 (
            .O(N__30483),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__6768 (
            .O(N__30480),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__6767 (
            .O(N__30477),
            .I(M_this_state_qZ0Z_10));
    InMux I__6766 (
            .O(N__30466),
            .I(N__30463));
    LocalMux I__6765 (
            .O(N__30463),
            .I(M_this_state_q_RNIR71EZ0Z_10));
    CascadeMux I__6764 (
            .O(N__30460),
            .I(N__30457));
    InMux I__6763 (
            .O(N__30457),
            .I(N__30454));
    LocalMux I__6762 (
            .O(N__30454),
            .I(\this_ppu.hspr_cry_0_c_inv_RNI1203 ));
    InMux I__6761 (
            .O(N__30451),
            .I(N__30439));
    InMux I__6760 (
            .O(N__30450),
            .I(N__30436));
    InMux I__6759 (
            .O(N__30449),
            .I(N__30427));
    InMux I__6758 (
            .O(N__30448),
            .I(N__30427));
    InMux I__6757 (
            .O(N__30447),
            .I(N__30427));
    InMux I__6756 (
            .O(N__30446),
            .I(N__30427));
    InMux I__6755 (
            .O(N__30445),
            .I(N__30418));
    InMux I__6754 (
            .O(N__30444),
            .I(N__30418));
    InMux I__6753 (
            .O(N__30443),
            .I(N__30418));
    InMux I__6752 (
            .O(N__30442),
            .I(N__30418));
    LocalMux I__6751 (
            .O(N__30439),
            .I(N__30409));
    LocalMux I__6750 (
            .O(N__30436),
            .I(N__30406));
    LocalMux I__6749 (
            .O(N__30427),
            .I(N__30401));
    LocalMux I__6748 (
            .O(N__30418),
            .I(N__30401));
    InMux I__6747 (
            .O(N__30417),
            .I(N__30396));
    InMux I__6746 (
            .O(N__30416),
            .I(N__30396));
    InMux I__6745 (
            .O(N__30415),
            .I(N__30387));
    InMux I__6744 (
            .O(N__30414),
            .I(N__30387));
    InMux I__6743 (
            .O(N__30413),
            .I(N__30387));
    InMux I__6742 (
            .O(N__30412),
            .I(N__30387));
    Odrv12 I__6741 (
            .O(N__30409),
            .I(N_332_0));
    Odrv4 I__6740 (
            .O(N__30406),
            .I(N_332_0));
    Odrv4 I__6739 (
            .O(N__30401),
            .I(N_332_0));
    LocalMux I__6738 (
            .O(N__30396),
            .I(N_332_0));
    LocalMux I__6737 (
            .O(N__30387),
            .I(N_332_0));
    CascadeMux I__6736 (
            .O(N__30376),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_ ));
    InMux I__6735 (
            .O(N__30373),
            .I(N__30370));
    LocalMux I__6734 (
            .O(N__30370),
            .I(\this_ppu.N_405 ));
    CascadeMux I__6733 (
            .O(N__30367),
            .I(N__30361));
    InMux I__6732 (
            .O(N__30366),
            .I(N__30356));
    InMux I__6731 (
            .O(N__30365),
            .I(N__30351));
    InMux I__6730 (
            .O(N__30364),
            .I(N__30351));
    InMux I__6729 (
            .O(N__30361),
            .I(N__30344));
    InMux I__6728 (
            .O(N__30360),
            .I(N__30344));
    InMux I__6727 (
            .O(N__30359),
            .I(N__30344));
    LocalMux I__6726 (
            .O(N__30356),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6725 (
            .O(N__30351),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__6724 (
            .O(N__30344),
            .I(M_this_state_qZ0Z_12));
    CascadeMux I__6723 (
            .O(N__30337),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_ ));
    CascadeMux I__6722 (
            .O(N__30334),
            .I(N__30331));
    InMux I__6721 (
            .O(N__30331),
            .I(N__30326));
    InMux I__6720 (
            .O(N__30330),
            .I(N__30323));
    InMux I__6719 (
            .O(N__30329),
            .I(N__30320));
    LocalMux I__6718 (
            .O(N__30326),
            .I(N__30315));
    LocalMux I__6717 (
            .O(N__30323),
            .I(N__30315));
    LocalMux I__6716 (
            .O(N__30320),
            .I(N__30310));
    Span4Mux_h I__6715 (
            .O(N__30315),
            .I(N__30310));
    Odrv4 I__6714 (
            .O(N__30310),
            .I(\this_ppu.N_324_0 ));
    CascadeMux I__6713 (
            .O(N__30307),
            .I(N__30304));
    CascadeBuf I__6712 (
            .O(N__30304),
            .I(N__30301));
    CascadeMux I__6711 (
            .O(N__30301),
            .I(N__30296));
    InMux I__6710 (
            .O(N__30300),
            .I(N__30293));
    CascadeMux I__6709 (
            .O(N__30299),
            .I(N__30290));
    InMux I__6708 (
            .O(N__30296),
            .I(N__30287));
    LocalMux I__6707 (
            .O(N__30293),
            .I(N__30283));
    InMux I__6706 (
            .O(N__30290),
            .I(N__30280));
    LocalMux I__6705 (
            .O(N__30287),
            .I(N__30277));
    InMux I__6704 (
            .O(N__30286),
            .I(N__30274));
    Span4Mux_h I__6703 (
            .O(N__30283),
            .I(N__30271));
    LocalMux I__6702 (
            .O(N__30280),
            .I(N__30266));
    Span4Mux_h I__6701 (
            .O(N__30277),
            .I(N__30266));
    LocalMux I__6700 (
            .O(N__30274),
            .I(\this_ppu.M_oamidx_qZ0Z_1 ));
    Odrv4 I__6699 (
            .O(N__30271),
            .I(\this_ppu.M_oamidx_qZ0Z_1 ));
    Odrv4 I__6698 (
            .O(N__30266),
            .I(\this_ppu.M_oamidx_qZ0Z_1 ));
    CascadeMux I__6697 (
            .O(N__30259),
            .I(N__30256));
    InMux I__6696 (
            .O(N__30256),
            .I(N__30253));
    LocalMux I__6695 (
            .O(N__30253),
            .I(N__30250));
    Odrv12 I__6694 (
            .O(N__30250),
            .I(\this_ppu.un1_M_oamidx_q_cry_0_THRU_CO ));
    InMux I__6693 (
            .O(N__30247),
            .I(\this_ppu.un1_M_oamidx_q_cry_0 ));
    CascadeMux I__6692 (
            .O(N__30244),
            .I(N__30241));
    InMux I__6691 (
            .O(N__30241),
            .I(N__30238));
    LocalMux I__6690 (
            .O(N__30238),
            .I(\this_ppu.un1_M_oamidx_q_cry_1_THRU_CO ));
    InMux I__6689 (
            .O(N__30235),
            .I(\this_ppu.un1_M_oamidx_q_cry_1 ));
    InMux I__6688 (
            .O(N__30232),
            .I(\this_ppu.un1_M_oamidx_q_cry_2 ));
    CascadeMux I__6687 (
            .O(N__30229),
            .I(N__30226));
    CascadeBuf I__6686 (
            .O(N__30226),
            .I(N__30223));
    CascadeMux I__6685 (
            .O(N__30223),
            .I(N__30220));
    InMux I__6684 (
            .O(N__30220),
            .I(N__30214));
    InMux I__6683 (
            .O(N__30219),
            .I(N__30211));
    InMux I__6682 (
            .O(N__30218),
            .I(N__30206));
    InMux I__6681 (
            .O(N__30217),
            .I(N__30206));
    LocalMux I__6680 (
            .O(N__30214),
            .I(N__30203));
    LocalMux I__6679 (
            .O(N__30211),
            .I(\this_ppu.M_oamidx_qZ1Z_2 ));
    LocalMux I__6678 (
            .O(N__30206),
            .I(\this_ppu.M_oamidx_qZ1Z_2 ));
    Odrv12 I__6677 (
            .O(N__30203),
            .I(\this_ppu.M_oamidx_qZ1Z_2 ));
    CascadeMux I__6676 (
            .O(N__30196),
            .I(N__30193));
    CascadeBuf I__6675 (
            .O(N__30193),
            .I(N__30190));
    CascadeMux I__6674 (
            .O(N__30190),
            .I(N__30187));
    InMux I__6673 (
            .O(N__30187),
            .I(N__30184));
    LocalMux I__6672 (
            .O(N__30184),
            .I(N__30179));
    CascadeMux I__6671 (
            .O(N__30183),
            .I(N__30175));
    InMux I__6670 (
            .O(N__30182),
            .I(N__30172));
    Span4Mux_v I__6669 (
            .O(N__30179),
            .I(N__30169));
    InMux I__6668 (
            .O(N__30178),
            .I(N__30165));
    InMux I__6667 (
            .O(N__30175),
            .I(N__30160));
    LocalMux I__6666 (
            .O(N__30172),
            .I(N__30155));
    Span4Mux_h I__6665 (
            .O(N__30169),
            .I(N__30155));
    InMux I__6664 (
            .O(N__30168),
            .I(N__30152));
    LocalMux I__6663 (
            .O(N__30165),
            .I(N__30149));
    InMux I__6662 (
            .O(N__30164),
            .I(N__30146));
    InMux I__6661 (
            .O(N__30163),
            .I(N__30143));
    LocalMux I__6660 (
            .O(N__30160),
            .I(N__30138));
    Span4Mux_h I__6659 (
            .O(N__30155),
            .I(N__30138));
    LocalMux I__6658 (
            .O(N__30152),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__6657 (
            .O(N__30149),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__6656 (
            .O(N__30146),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__6655 (
            .O(N__30143),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__6654 (
            .O(N__30138),
            .I(M_this_ppu_oam_addr_3));
    CascadeMux I__6653 (
            .O(N__30127),
            .I(N__30124));
    CascadeBuf I__6652 (
            .O(N__30124),
            .I(N__30121));
    CascadeMux I__6651 (
            .O(N__30121),
            .I(N__30116));
    CascadeMux I__6650 (
            .O(N__30120),
            .I(N__30113));
    CascadeMux I__6649 (
            .O(N__30119),
            .I(N__30110));
    InMux I__6648 (
            .O(N__30116),
            .I(N__30107));
    InMux I__6647 (
            .O(N__30113),
            .I(N__30102));
    InMux I__6646 (
            .O(N__30110),
            .I(N__30102));
    LocalMux I__6645 (
            .O(N__30107),
            .I(N__30099));
    LocalMux I__6644 (
            .O(N__30102),
            .I(N__30094));
    Span4Mux_h I__6643 (
            .O(N__30099),
            .I(N__30094));
    Odrv4 I__6642 (
            .O(N__30094),
            .I(\this_ppu.M_oamidx_qZ0Z_3 ));
    CascadeMux I__6641 (
            .O(N__30091),
            .I(N__30088));
    CascadeBuf I__6640 (
            .O(N__30088),
            .I(N__30085));
    CascadeMux I__6639 (
            .O(N__30085),
            .I(N__30082));
    InMux I__6638 (
            .O(N__30082),
            .I(N__30078));
    InMux I__6637 (
            .O(N__30081),
            .I(N__30074));
    LocalMux I__6636 (
            .O(N__30078),
            .I(N__30071));
    CascadeMux I__6635 (
            .O(N__30077),
            .I(N__30067));
    LocalMux I__6634 (
            .O(N__30074),
            .I(N__30063));
    Span4Mux_v I__6633 (
            .O(N__30071),
            .I(N__30060));
    InMux I__6632 (
            .O(N__30070),
            .I(N__30057));
    InMux I__6631 (
            .O(N__30067),
            .I(N__30054));
    InMux I__6630 (
            .O(N__30066),
            .I(N__30051));
    Span4Mux_v I__6629 (
            .O(N__30063),
            .I(N__30046));
    Span4Mux_h I__6628 (
            .O(N__30060),
            .I(N__30046));
    LocalMux I__6627 (
            .O(N__30057),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__6626 (
            .O(N__30054),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__6625 (
            .O(N__30051),
            .I(M_this_ppu_oam_addr_2));
    Odrv4 I__6624 (
            .O(N__30046),
            .I(M_this_ppu_oam_addr_2));
    InMux I__6623 (
            .O(N__30037),
            .I(N__30034));
    LocalMux I__6622 (
            .O(N__30034),
            .I(N__30031));
    Span4Mux_h I__6621 (
            .O(N__30031),
            .I(N__30028));
    Odrv4 I__6620 (
            .O(N__30028),
            .I(\this_ppu.M_state_q_srsts_0_a3_0_o2_0_6 ));
    InMux I__6619 (
            .O(N__30025),
            .I(N__30016));
    InMux I__6618 (
            .O(N__30024),
            .I(N__30011));
    InMux I__6617 (
            .O(N__30023),
            .I(N__30011));
    CascadeMux I__6616 (
            .O(N__30022),
            .I(N__30007));
    InMux I__6615 (
            .O(N__30021),
            .I(N__30004));
    InMux I__6614 (
            .O(N__30020),
            .I(N__30001));
    InMux I__6613 (
            .O(N__30019),
            .I(N__29995));
    LocalMux I__6612 (
            .O(N__30016),
            .I(N__29990));
    LocalMux I__6611 (
            .O(N__30011),
            .I(N__29990));
    InMux I__6610 (
            .O(N__30010),
            .I(N__29987));
    InMux I__6609 (
            .O(N__30007),
            .I(N__29984));
    LocalMux I__6608 (
            .O(N__30004),
            .I(N__29977));
    LocalMux I__6607 (
            .O(N__30001),
            .I(N__29977));
    InMux I__6606 (
            .O(N__30000),
            .I(N__29974));
    InMux I__6605 (
            .O(N__29999),
            .I(N__29969));
    InMux I__6604 (
            .O(N__29998),
            .I(N__29969));
    LocalMux I__6603 (
            .O(N__29995),
            .I(N__29965));
    Span4Mux_v I__6602 (
            .O(N__29990),
            .I(N__29962));
    LocalMux I__6601 (
            .O(N__29987),
            .I(N__29957));
    LocalMux I__6600 (
            .O(N__29984),
            .I(N__29957));
    InMux I__6599 (
            .O(N__29983),
            .I(N__29954));
    InMux I__6598 (
            .O(N__29982),
            .I(N__29951));
    Span4Mux_v I__6597 (
            .O(N__29977),
            .I(N__29944));
    LocalMux I__6596 (
            .O(N__29974),
            .I(N__29944));
    LocalMux I__6595 (
            .O(N__29969),
            .I(N__29944));
    InMux I__6594 (
            .O(N__29968),
            .I(N__29941));
    Span4Mux_v I__6593 (
            .O(N__29965),
            .I(N__29938));
    Span4Mux_h I__6592 (
            .O(N__29962),
            .I(N__29931));
    Span4Mux_h I__6591 (
            .O(N__29957),
            .I(N__29931));
    LocalMux I__6590 (
            .O(N__29954),
            .I(N__29931));
    LocalMux I__6589 (
            .O(N__29951),
            .I(N__29928));
    Span4Mux_v I__6588 (
            .O(N__29944),
            .I(N__29925));
    LocalMux I__6587 (
            .O(N__29941),
            .I(N__29922));
    Span4Mux_h I__6586 (
            .O(N__29938),
            .I(N__29917));
    Span4Mux_v I__6585 (
            .O(N__29931),
            .I(N__29917));
    Span4Mux_h I__6584 (
            .O(N__29928),
            .I(N__29914));
    Span4Mux_h I__6583 (
            .O(N__29925),
            .I(N__29911));
    Span4Mux_v I__6582 (
            .O(N__29922),
            .I(N__29906));
    Span4Mux_h I__6581 (
            .O(N__29917),
            .I(N__29906));
    Span4Mux_v I__6580 (
            .O(N__29914),
            .I(N__29901));
    Span4Mux_v I__6579 (
            .O(N__29911),
            .I(N__29901));
    Odrv4 I__6578 (
            .O(N__29906),
            .I(\this_ppu.N_228_0_i_1_0 ));
    Odrv4 I__6577 (
            .O(N__29901),
            .I(\this_ppu.N_228_0_i_1_0 ));
    CascadeMux I__6576 (
            .O(N__29896),
            .I(N__29893));
    CascadeBuf I__6575 (
            .O(N__29893),
            .I(N__29889));
    InMux I__6574 (
            .O(N__29892),
            .I(N__29886));
    CascadeMux I__6573 (
            .O(N__29889),
            .I(N__29881));
    LocalMux I__6572 (
            .O(N__29886),
            .I(N__29878));
    CascadeMux I__6571 (
            .O(N__29885),
            .I(N__29875));
    CascadeMux I__6570 (
            .O(N__29884),
            .I(N__29872));
    InMux I__6569 (
            .O(N__29881),
            .I(N__29869));
    Span4Mux_v I__6568 (
            .O(N__29878),
            .I(N__29866));
    InMux I__6567 (
            .O(N__29875),
            .I(N__29861));
    InMux I__6566 (
            .O(N__29872),
            .I(N__29861));
    LocalMux I__6565 (
            .O(N__29869),
            .I(N__29858));
    Odrv4 I__6564 (
            .O(N__29866),
            .I(\this_ppu.M_oamidx_qZ0Z_0 ));
    LocalMux I__6563 (
            .O(N__29861),
            .I(\this_ppu.M_oamidx_qZ0Z_0 ));
    Odrv12 I__6562 (
            .O(N__29858),
            .I(\this_ppu.M_oamidx_qZ0Z_0 ));
    InMux I__6561 (
            .O(N__29851),
            .I(N__29848));
    LocalMux I__6560 (
            .O(N__29848),
            .I(N__29844));
    InMux I__6559 (
            .O(N__29847),
            .I(N__29840));
    Span4Mux_h I__6558 (
            .O(N__29844),
            .I(N__29837));
    InMux I__6557 (
            .O(N__29843),
            .I(N__29834));
    LocalMux I__6556 (
            .O(N__29840),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv4 I__6555 (
            .O(N__29837),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    LocalMux I__6554 (
            .O(N__29834),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    InMux I__6553 (
            .O(N__29827),
            .I(N__29824));
    LocalMux I__6552 (
            .O(N__29824),
            .I(\this_ppu.N_255 ));
    InMux I__6551 (
            .O(N__29821),
            .I(N__29817));
    InMux I__6550 (
            .O(N__29820),
            .I(N__29814));
    LocalMux I__6549 (
            .O(N__29817),
            .I(N__29810));
    LocalMux I__6548 (
            .O(N__29814),
            .I(N__29807));
    InMux I__6547 (
            .O(N__29813),
            .I(N__29804));
    Odrv4 I__6546 (
            .O(N__29810),
            .I(\this_ppu.N_756_0 ));
    Odrv4 I__6545 (
            .O(N__29807),
            .I(\this_ppu.N_756_0 ));
    LocalMux I__6544 (
            .O(N__29804),
            .I(\this_ppu.N_756_0 ));
    InMux I__6543 (
            .O(N__29797),
            .I(N__29791));
    InMux I__6542 (
            .O(N__29796),
            .I(N__29791));
    LocalMux I__6541 (
            .O(N__29791),
            .I(\this_ppu.un1_M_vaddress_q_c2 ));
    InMux I__6540 (
            .O(N__29788),
            .I(N__29779));
    InMux I__6539 (
            .O(N__29787),
            .I(N__29779));
    InMux I__6538 (
            .O(N__29786),
            .I(N__29779));
    LocalMux I__6537 (
            .O(N__29779),
            .I(\this_ppu.un1_M_vaddress_q_c5 ));
    SRMux I__6536 (
            .O(N__29776),
            .I(N__29773));
    LocalMux I__6535 (
            .O(N__29773),
            .I(N__29770));
    Span4Mux_v I__6534 (
            .O(N__29770),
            .I(N__29766));
    SRMux I__6533 (
            .O(N__29769),
            .I(N__29763));
    Span4Mux_h I__6532 (
            .O(N__29766),
            .I(N__29760));
    LocalMux I__6531 (
            .O(N__29763),
            .I(N__29757));
    Span4Mux_h I__6530 (
            .O(N__29760),
            .I(N__29751));
    Span4Mux_v I__6529 (
            .O(N__29757),
            .I(N__29751));
    SRMux I__6528 (
            .O(N__29756),
            .I(N__29748));
    Sp12to4 I__6527 (
            .O(N__29751),
            .I(N__29745));
    LocalMux I__6526 (
            .O(N__29748),
            .I(N__29742));
    Odrv12 I__6525 (
            .O(N__29745),
            .I(\this_ppu.M_last_q_RNIITCPC ));
    Odrv4 I__6524 (
            .O(N__29742),
            .I(\this_ppu.M_last_q_RNIITCPC ));
    InMux I__6523 (
            .O(N__29737),
            .I(\this_ppu.un1_M_oam_cache_read_data_2_cry_8 ));
    InMux I__6522 (
            .O(N__29734),
            .I(N__29731));
    LocalMux I__6521 (
            .O(N__29731),
            .I(N__29726));
    InMux I__6520 (
            .O(N__29730),
            .I(N__29723));
    InMux I__6519 (
            .O(N__29729),
            .I(N__29720));
    Span4Mux_h I__6518 (
            .O(N__29726),
            .I(N__29715));
    LocalMux I__6517 (
            .O(N__29723),
            .I(N__29715));
    LocalMux I__6516 (
            .O(N__29720),
            .I(N__29712));
    Odrv4 I__6515 (
            .O(N__29715),
            .I(\this_ppu.N_242_0 ));
    Odrv4 I__6514 (
            .O(N__29712),
            .I(\this_ppu.N_242_0 ));
    InMux I__6513 (
            .O(N__29707),
            .I(N__29704));
    LocalMux I__6512 (
            .O(N__29704),
            .I(N__29701));
    Span4Mux_v I__6511 (
            .O(N__29701),
            .I(N__29698));
    Span4Mux_h I__6510 (
            .O(N__29698),
            .I(N__29695));
    Odrv4 I__6509 (
            .O(N__29695),
            .I(\this_ppu.oam_cache.mem_4 ));
    InMux I__6508 (
            .O(N__29692),
            .I(N__29689));
    LocalMux I__6507 (
            .O(N__29689),
            .I(N__29686));
    Odrv12 I__6506 (
            .O(N__29686),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_4 ));
    InMux I__6505 (
            .O(N__29683),
            .I(N__29679));
    InMux I__6504 (
            .O(N__29682),
            .I(N__29676));
    LocalMux I__6503 (
            .O(N__29679),
            .I(N__29671));
    LocalMux I__6502 (
            .O(N__29676),
            .I(N__29667));
    InMux I__6501 (
            .O(N__29675),
            .I(N__29664));
    InMux I__6500 (
            .O(N__29674),
            .I(N__29661));
    Span4Mux_h I__6499 (
            .O(N__29671),
            .I(N__29658));
    InMux I__6498 (
            .O(N__29670),
            .I(N__29655));
    Span4Mux_v I__6497 (
            .O(N__29667),
            .I(N__29650));
    LocalMux I__6496 (
            .O(N__29664),
            .I(N__29650));
    LocalMux I__6495 (
            .O(N__29661),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_7 ));
    Odrv4 I__6494 (
            .O(N__29658),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_7 ));
    LocalMux I__6493 (
            .O(N__29655),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_7 ));
    Odrv4 I__6492 (
            .O(N__29650),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_7 ));
    InMux I__6491 (
            .O(N__29641),
            .I(N__29637));
    InMux I__6490 (
            .O(N__29640),
            .I(N__29634));
    LocalMux I__6489 (
            .O(N__29637),
            .I(N__29629));
    LocalMux I__6488 (
            .O(N__29634),
            .I(N__29626));
    InMux I__6487 (
            .O(N__29633),
            .I(N__29622));
    InMux I__6486 (
            .O(N__29632),
            .I(N__29619));
    Span4Mux_h I__6485 (
            .O(N__29629),
            .I(N__29614));
    Span4Mux_v I__6484 (
            .O(N__29626),
            .I(N__29614));
    InMux I__6483 (
            .O(N__29625),
            .I(N__29611));
    LocalMux I__6482 (
            .O(N__29622),
            .I(N__29608));
    LocalMux I__6481 (
            .O(N__29619),
            .I(N__29605));
    Span4Mux_v I__6480 (
            .O(N__29614),
            .I(N__29602));
    LocalMux I__6479 (
            .O(N__29611),
            .I(N__29599));
    Span12Mux_v I__6478 (
            .O(N__29608),
            .I(N__29596));
    Sp12to4 I__6477 (
            .O(N__29605),
            .I(N__29593));
    Span4Mux_v I__6476 (
            .O(N__29602),
            .I(N__29588));
    Span4Mux_v I__6475 (
            .O(N__29599),
            .I(N__29588));
    Odrv12 I__6474 (
            .O(N__29596),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv12 I__6473 (
            .O(N__29593),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv4 I__6472 (
            .O(N__29588),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    InMux I__6471 (
            .O(N__29581),
            .I(N__29576));
    InMux I__6470 (
            .O(N__29580),
            .I(N__29573));
    InMux I__6469 (
            .O(N__29579),
            .I(N__29570));
    LocalMux I__6468 (
            .O(N__29576),
            .I(N__29567));
    LocalMux I__6467 (
            .O(N__29573),
            .I(N__29564));
    LocalMux I__6466 (
            .O(N__29570),
            .I(N__29561));
    Span12Mux_h I__6465 (
            .O(N__29567),
            .I(N__29557));
    Span12Mux_v I__6464 (
            .O(N__29564),
            .I(N__29553));
    Span4Mux_h I__6463 (
            .O(N__29561),
            .I(N__29550));
    InMux I__6462 (
            .O(N__29560),
            .I(N__29547));
    Span12Mux_v I__6461 (
            .O(N__29557),
            .I(N__29544));
    InMux I__6460 (
            .O(N__29556),
            .I(N__29541));
    Odrv12 I__6459 (
            .O(N__29553),
            .I(\this_ppu.N_772_0 ));
    Odrv4 I__6458 (
            .O(N__29550),
            .I(\this_ppu.N_772_0 ));
    LocalMux I__6457 (
            .O(N__29547),
            .I(\this_ppu.N_772_0 ));
    Odrv12 I__6456 (
            .O(N__29544),
            .I(\this_ppu.N_772_0 ));
    LocalMux I__6455 (
            .O(N__29541),
            .I(\this_ppu.N_772_0 ));
    InMux I__6454 (
            .O(N__29530),
            .I(N__29527));
    LocalMux I__6453 (
            .O(N__29527),
            .I(N__29524));
    Odrv12 I__6452 (
            .O(N__29524),
            .I(\this_ppu.N_760_0 ));
    InMux I__6451 (
            .O(N__29521),
            .I(N__29515));
    InMux I__6450 (
            .O(N__29520),
            .I(N__29511));
    InMux I__6449 (
            .O(N__29519),
            .I(N__29506));
    InMux I__6448 (
            .O(N__29518),
            .I(N__29506));
    LocalMux I__6447 (
            .O(N__29515),
            .I(N__29503));
    InMux I__6446 (
            .O(N__29514),
            .I(N__29500));
    LocalMux I__6445 (
            .O(N__29511),
            .I(N__29497));
    LocalMux I__6444 (
            .O(N__29506),
            .I(N__29494));
    Span4Mux_v I__6443 (
            .O(N__29503),
            .I(N__29489));
    LocalMux I__6442 (
            .O(N__29500),
            .I(N__29489));
    Span4Mux_v I__6441 (
            .O(N__29497),
            .I(N__29486));
    Odrv12 I__6440 (
            .O(N__29494),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__6439 (
            .O(N__29489),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    Odrv4 I__6438 (
            .O(N__29486),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    CascadeMux I__6437 (
            .O(N__29479),
            .I(\this_ppu.N_799_cascade_ ));
    InMux I__6436 (
            .O(N__29476),
            .I(N__29471));
    InMux I__6435 (
            .O(N__29475),
            .I(N__29468));
    InMux I__6434 (
            .O(N__29474),
            .I(N__29465));
    LocalMux I__6433 (
            .O(N__29471),
            .I(N__29462));
    LocalMux I__6432 (
            .O(N__29468),
            .I(\this_ppu.N_779_0 ));
    LocalMux I__6431 (
            .O(N__29465),
            .I(\this_ppu.N_779_0 ));
    Odrv4 I__6430 (
            .O(N__29462),
            .I(\this_ppu.N_779_0 ));
    CascadeMux I__6429 (
            .O(N__29455),
            .I(N__29452));
    InMux I__6428 (
            .O(N__29452),
            .I(N__29444));
    CascadeMux I__6427 (
            .O(N__29451),
            .I(N__29440));
    InMux I__6426 (
            .O(N__29450),
            .I(N__29437));
    InMux I__6425 (
            .O(N__29449),
            .I(N__29433));
    InMux I__6424 (
            .O(N__29448),
            .I(N__29430));
    CascadeMux I__6423 (
            .O(N__29447),
            .I(N__29427));
    LocalMux I__6422 (
            .O(N__29444),
            .I(N__29424));
    InMux I__6421 (
            .O(N__29443),
            .I(N__29419));
    InMux I__6420 (
            .O(N__29440),
            .I(N__29419));
    LocalMux I__6419 (
            .O(N__29437),
            .I(N__29416));
    CascadeMux I__6418 (
            .O(N__29436),
            .I(N__29412));
    LocalMux I__6417 (
            .O(N__29433),
            .I(N__29407));
    LocalMux I__6416 (
            .O(N__29430),
            .I(N__29407));
    InMux I__6415 (
            .O(N__29427),
            .I(N__29404));
    Span4Mux_v I__6414 (
            .O(N__29424),
            .I(N__29399));
    LocalMux I__6413 (
            .O(N__29419),
            .I(N__29399));
    Span4Mux_v I__6412 (
            .O(N__29416),
            .I(N__29396));
    InMux I__6411 (
            .O(N__29415),
            .I(N__29393));
    InMux I__6410 (
            .O(N__29412),
            .I(N__29390));
    Span4Mux_v I__6409 (
            .O(N__29407),
            .I(N__29385));
    LocalMux I__6408 (
            .O(N__29404),
            .I(N__29385));
    Span4Mux_v I__6407 (
            .O(N__29399),
            .I(N__29380));
    Span4Mux_h I__6406 (
            .O(N__29396),
            .I(N__29380));
    LocalMux I__6405 (
            .O(N__29393),
            .I(N__29377));
    LocalMux I__6404 (
            .O(N__29390),
            .I(N__29374));
    Span4Mux_h I__6403 (
            .O(N__29385),
            .I(N__29371));
    Odrv4 I__6402 (
            .O(N__29380),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__6401 (
            .O(N__29377),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__6400 (
            .O(N__29374),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__6399 (
            .O(N__29371),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    InMux I__6398 (
            .O(N__29362),
            .I(N__29359));
    LocalMux I__6397 (
            .O(N__29359),
            .I(\this_ppu.N_267 ));
    CascadeMux I__6396 (
            .O(N__29356),
            .I(N__29353));
    InMux I__6395 (
            .O(N__29353),
            .I(N__29349));
    InMux I__6394 (
            .O(N__29352),
            .I(N__29346));
    LocalMux I__6393 (
            .O(N__29349),
            .I(N__29342));
    LocalMux I__6392 (
            .O(N__29346),
            .I(N__29339));
    InMux I__6391 (
            .O(N__29345),
            .I(N__29334));
    Span4Mux_h I__6390 (
            .O(N__29342),
            .I(N__29331));
    Span4Mux_v I__6389 (
            .O(N__29339),
            .I(N__29327));
    CascadeMux I__6388 (
            .O(N__29338),
            .I(N__29324));
    CascadeMux I__6387 (
            .O(N__29337),
            .I(N__29320));
    LocalMux I__6386 (
            .O(N__29334),
            .I(N__29316));
    Span4Mux_v I__6385 (
            .O(N__29331),
            .I(N__29313));
    InMux I__6384 (
            .O(N__29330),
            .I(N__29310));
    Span4Mux_h I__6383 (
            .O(N__29327),
            .I(N__29307));
    InMux I__6382 (
            .O(N__29324),
            .I(N__29300));
    InMux I__6381 (
            .O(N__29323),
            .I(N__29300));
    InMux I__6380 (
            .O(N__29320),
            .I(N__29300));
    InMux I__6379 (
            .O(N__29319),
            .I(N__29297));
    Span12Mux_h I__6378 (
            .O(N__29316),
            .I(N__29294));
    Span4Mux_h I__6377 (
            .O(N__29313),
            .I(N__29289));
    LocalMux I__6376 (
            .O(N__29310),
            .I(N__29289));
    Odrv4 I__6375 (
            .O(N__29307),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__6374 (
            .O(N__29300),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__6373 (
            .O(N__29297),
            .I(M_this_ppu_vram_addr_0));
    Odrv12 I__6372 (
            .O(N__29294),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__6371 (
            .O(N__29289),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__6370 (
            .O(N__29278),
            .I(N__29275));
    InMux I__6369 (
            .O(N__29275),
            .I(N__29272));
    LocalMux I__6368 (
            .O(N__29272),
            .I(N__29268));
    CascadeMux I__6367 (
            .O(N__29271),
            .I(N__29265));
    Span4Mux_h I__6366 (
            .O(N__29268),
            .I(N__29262));
    InMux I__6365 (
            .O(N__29265),
            .I(N__29259));
    Odrv4 I__6364 (
            .O(N__29262),
            .I(M_this_scroll_qZ0Z_8));
    LocalMux I__6363 (
            .O(N__29259),
            .I(M_this_scroll_qZ0Z_8));
    InMux I__6362 (
            .O(N__29254),
            .I(N__29251));
    LocalMux I__6361 (
            .O(N__29251),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12 ));
    InMux I__6360 (
            .O(N__29248),
            .I(N__29245));
    LocalMux I__6359 (
            .O(N__29245),
            .I(dma_axb3));
    CascadeMux I__6358 (
            .O(N__29242),
            .I(this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_));
    IoInMux I__6357 (
            .O(N__29239),
            .I(N__29236));
    LocalMux I__6356 (
            .O(N__29236),
            .I(N__29233));
    IoSpan4Mux I__6355 (
            .O(N__29233),
            .I(N__29230));
    Span4Mux_s2_h I__6354 (
            .O(N__29230),
            .I(N__29226));
    InMux I__6353 (
            .O(N__29229),
            .I(N__29220));
    Span4Mux_h I__6352 (
            .O(N__29226),
            .I(N__29217));
    InMux I__6351 (
            .O(N__29225),
            .I(N__29214));
    CascadeMux I__6350 (
            .O(N__29224),
            .I(N__29211));
    InMux I__6349 (
            .O(N__29223),
            .I(N__29208));
    LocalMux I__6348 (
            .O(N__29220),
            .I(N__29205));
    Span4Mux_h I__6347 (
            .O(N__29217),
            .I(N__29200));
    LocalMux I__6346 (
            .O(N__29214),
            .I(N__29200));
    InMux I__6345 (
            .O(N__29211),
            .I(N__29197));
    LocalMux I__6344 (
            .O(N__29208),
            .I(N__29194));
    Span4Mux_v I__6343 (
            .O(N__29205),
            .I(N__29191));
    Span4Mux_v I__6342 (
            .O(N__29200),
            .I(N__29186));
    LocalMux I__6341 (
            .O(N__29197),
            .I(N__29186));
    Span4Mux_v I__6340 (
            .O(N__29194),
            .I(N__29183));
    Span4Mux_h I__6339 (
            .O(N__29191),
            .I(N__29180));
    Span4Mux_h I__6338 (
            .O(N__29186),
            .I(N__29177));
    Sp12to4 I__6337 (
            .O(N__29183),
            .I(N__29174));
    Span4Mux_h I__6336 (
            .O(N__29180),
            .I(N__29169));
    Span4Mux_v I__6335 (
            .O(N__29177),
            .I(N__29169));
    Span12Mux_s9_h I__6334 (
            .O(N__29174),
            .I(N__29166));
    Span4Mux_h I__6333 (
            .O(N__29169),
            .I(N__29163));
    Odrv12 I__6332 (
            .O(N__29166),
            .I(dma_0));
    Odrv4 I__6331 (
            .O(N__29163),
            .I(dma_0));
    InMux I__6330 (
            .O(N__29158),
            .I(N__29155));
    LocalMux I__6329 (
            .O(N__29155),
            .I(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10 ));
    CascadeMux I__6328 (
            .O(N__29152),
            .I(\this_ppu.N_414_1_cascade_ ));
    CascadeMux I__6327 (
            .O(N__29149),
            .I(N__29145));
    InMux I__6326 (
            .O(N__29148),
            .I(N__29142));
    InMux I__6325 (
            .O(N__29145),
            .I(N__29136));
    LocalMux I__6324 (
            .O(N__29142),
            .I(N__29133));
    InMux I__6323 (
            .O(N__29141),
            .I(N__29130));
    CascadeMux I__6322 (
            .O(N__29140),
            .I(N__29127));
    InMux I__6321 (
            .O(N__29139),
            .I(N__29124));
    LocalMux I__6320 (
            .O(N__29136),
            .I(N__29121));
    Span4Mux_v I__6319 (
            .O(N__29133),
            .I(N__29116));
    LocalMux I__6318 (
            .O(N__29130),
            .I(N__29116));
    InMux I__6317 (
            .O(N__29127),
            .I(N__29112));
    LocalMux I__6316 (
            .O(N__29124),
            .I(N__29109));
    Span4Mux_v I__6315 (
            .O(N__29121),
            .I(N__29106));
    Span4Mux_v I__6314 (
            .O(N__29116),
            .I(N__29103));
    InMux I__6313 (
            .O(N__29115),
            .I(N__29100));
    LocalMux I__6312 (
            .O(N__29112),
            .I(N__29095));
    Span12Mux_v I__6311 (
            .O(N__29109),
            .I(N__29095));
    Span4Mux_h I__6310 (
            .O(N__29106),
            .I(N__29090));
    Span4Mux_h I__6309 (
            .O(N__29103),
            .I(N__29090));
    LocalMux I__6308 (
            .O(N__29100),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv12 I__6307 (
            .O(N__29095),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__6306 (
            .O(N__29090),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    InMux I__6305 (
            .O(N__29083),
            .I(N__29080));
    LocalMux I__6304 (
            .O(N__29080),
            .I(N__29077));
    Odrv4 I__6303 (
            .O(N__29077),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__6302 (
            .O(N__29074),
            .I(N__29071));
    LocalMux I__6301 (
            .O(N__29071),
            .I(N__29068));
    Odrv12 I__6300 (
            .O(N__29068),
            .I(M_this_oam_ram_write_data_9));
    CEMux I__6299 (
            .O(N__29065),
            .I(N__29061));
    CEMux I__6298 (
            .O(N__29064),
            .I(N__29058));
    LocalMux I__6297 (
            .O(N__29061),
            .I(N__29054));
    LocalMux I__6296 (
            .O(N__29058),
            .I(N__29050));
    CEMux I__6295 (
            .O(N__29057),
            .I(N__29047));
    Span4Mux_h I__6294 (
            .O(N__29054),
            .I(N__29043));
    CEMux I__6293 (
            .O(N__29053),
            .I(N__29040));
    Span4Mux_v I__6292 (
            .O(N__29050),
            .I(N__29036));
    LocalMux I__6291 (
            .O(N__29047),
            .I(N__29033));
    CEMux I__6290 (
            .O(N__29046),
            .I(N__29030));
    Span4Mux_h I__6289 (
            .O(N__29043),
            .I(N__29025));
    LocalMux I__6288 (
            .O(N__29040),
            .I(N__29025));
    CEMux I__6287 (
            .O(N__29039),
            .I(N__29022));
    Span4Mux_h I__6286 (
            .O(N__29036),
            .I(N__29015));
    Span4Mux_v I__6285 (
            .O(N__29033),
            .I(N__29015));
    LocalMux I__6284 (
            .O(N__29030),
            .I(N__29015));
    Span4Mux_v I__6283 (
            .O(N__29025),
            .I(N__29010));
    LocalMux I__6282 (
            .O(N__29022),
            .I(N__29010));
    Odrv4 I__6281 (
            .O(N__29015),
            .I(N_1294_0));
    Odrv4 I__6280 (
            .O(N__29010),
            .I(N_1294_0));
    InMux I__6279 (
            .O(N__29005),
            .I(N__29002));
    LocalMux I__6278 (
            .O(N__29002),
            .I(N__28999));
    Odrv12 I__6277 (
            .O(N__28999),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__6276 (
            .O(N__28996),
            .I(N__28993));
    LocalMux I__6275 (
            .O(N__28993),
            .I(N__28990));
    Span4Mux_v I__6274 (
            .O(N__28990),
            .I(N__28987));
    Span4Mux_h I__6273 (
            .O(N__28987),
            .I(N__28984));
    Odrv4 I__6272 (
            .O(N__28984),
            .I(M_this_oam_ram_write_data_14));
    InMux I__6271 (
            .O(N__28981),
            .I(N__28978));
    LocalMux I__6270 (
            .O(N__28978),
            .I(N__28975));
    Span12Mux_v I__6269 (
            .O(N__28975),
            .I(N__28972));
    Odrv12 I__6268 (
            .O(N__28972),
            .I(\this_ppu.oam_cache.mem_6 ));
    InMux I__6267 (
            .O(N__28969),
            .I(N__28966));
    LocalMux I__6266 (
            .O(N__28966),
            .I(N__28963));
    Odrv12 I__6265 (
            .O(N__28963),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_6 ));
    CascadeMux I__6264 (
            .O(N__28960),
            .I(\this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_ ));
    InMux I__6263 (
            .O(N__28957),
            .I(N__28951));
    InMux I__6262 (
            .O(N__28956),
            .I(N__28951));
    LocalMux I__6261 (
            .O(N__28951),
            .I(N__28944));
    InMux I__6260 (
            .O(N__28950),
            .I(N__28941));
    InMux I__6259 (
            .O(N__28949),
            .I(N__28938));
    InMux I__6258 (
            .O(N__28948),
            .I(N__28933));
    InMux I__6257 (
            .O(N__28947),
            .I(N__28933));
    Span4Mux_h I__6256 (
            .O(N__28944),
            .I(N__28930));
    LocalMux I__6255 (
            .O(N__28941),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__6254 (
            .O(N__28938),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__6253 (
            .O(N__28933),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__6252 (
            .O(N__28930),
            .I(M_this_state_qZ0Z_8));
    CascadeMux I__6251 (
            .O(N__28921),
            .I(N__28917));
    InMux I__6250 (
            .O(N__28920),
            .I(N__28914));
    InMux I__6249 (
            .O(N__28917),
            .I(N__28911));
    LocalMux I__6248 (
            .O(N__28914),
            .I(N_260));
    LocalMux I__6247 (
            .O(N__28911),
            .I(N_260));
    InMux I__6246 (
            .O(N__28906),
            .I(N__28903));
    LocalMux I__6245 (
            .O(N__28903),
            .I(\this_ppu.N_406 ));
    SRMux I__6244 (
            .O(N__28900),
            .I(N__28867));
    SRMux I__6243 (
            .O(N__28899),
            .I(N__28867));
    SRMux I__6242 (
            .O(N__28898),
            .I(N__28867));
    SRMux I__6241 (
            .O(N__28897),
            .I(N__28867));
    SRMux I__6240 (
            .O(N__28896),
            .I(N__28867));
    SRMux I__6239 (
            .O(N__28895),
            .I(N__28867));
    SRMux I__6238 (
            .O(N__28894),
            .I(N__28867));
    SRMux I__6237 (
            .O(N__28893),
            .I(N__28867));
    SRMux I__6236 (
            .O(N__28892),
            .I(N__28867));
    SRMux I__6235 (
            .O(N__28891),
            .I(N__28867));
    SRMux I__6234 (
            .O(N__28890),
            .I(N__28867));
    GlobalMux I__6233 (
            .O(N__28867),
            .I(N__28864));
    gio2CtrlBuf I__6232 (
            .O(N__28864),
            .I(N_504_g));
    CascadeMux I__6231 (
            .O(N__28861),
            .I(N__28858));
    CascadeBuf I__6230 (
            .O(N__28858),
            .I(N__28855));
    CascadeMux I__6229 (
            .O(N__28855),
            .I(N__28852));
    InMux I__6228 (
            .O(N__28852),
            .I(N__28849));
    LocalMux I__6227 (
            .O(N__28849),
            .I(N__28846));
    Odrv12 I__6226 (
            .O(N__28846),
            .I(\this_ppu.N_17_0 ));
    CascadeMux I__6225 (
            .O(N__28843),
            .I(\this_ppu.N_329_0_cascade_ ));
    InMux I__6224 (
            .O(N__28840),
            .I(N__28836));
    InMux I__6223 (
            .O(N__28839),
            .I(N__28833));
    LocalMux I__6222 (
            .O(N__28836),
            .I(\this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2 ));
    LocalMux I__6221 (
            .O(N__28833),
            .I(\this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2 ));
    CascadeMux I__6220 (
            .O(N__28828),
            .I(N__28825));
    CascadeBuf I__6219 (
            .O(N__28825),
            .I(N__28822));
    CascadeMux I__6218 (
            .O(N__28822),
            .I(N__28819));
    InMux I__6217 (
            .O(N__28819),
            .I(N__28816));
    LocalMux I__6216 (
            .O(N__28816),
            .I(N__28813));
    Span4Mux_h I__6215 (
            .O(N__28813),
            .I(N__28810));
    Odrv4 I__6214 (
            .O(N__28810),
            .I(\this_ppu.N_21_0 ));
    InMux I__6213 (
            .O(N__28807),
            .I(N__28801));
    InMux I__6212 (
            .O(N__28806),
            .I(N__28798));
    InMux I__6211 (
            .O(N__28805),
            .I(N__28795));
    InMux I__6210 (
            .O(N__28804),
            .I(N__28792));
    LocalMux I__6209 (
            .O(N__28801),
            .I(\this_ppu.un1_M_oamcurr_q_2_c3 ));
    LocalMux I__6208 (
            .O(N__28798),
            .I(\this_ppu.un1_M_oamcurr_q_2_c3 ));
    LocalMux I__6207 (
            .O(N__28795),
            .I(\this_ppu.un1_M_oamcurr_q_2_c3 ));
    LocalMux I__6206 (
            .O(N__28792),
            .I(\this_ppu.un1_M_oamcurr_q_2_c3 ));
    CascadeMux I__6205 (
            .O(N__28783),
            .I(N__28780));
    CascadeBuf I__6204 (
            .O(N__28780),
            .I(N__28777));
    CascadeMux I__6203 (
            .O(N__28777),
            .I(N__28774));
    InMux I__6202 (
            .O(N__28774),
            .I(N__28771));
    LocalMux I__6201 (
            .O(N__28771),
            .I(N__28768));
    Odrv12 I__6200 (
            .O(N__28768),
            .I(\this_ppu.N_23_0 ));
    InMux I__6199 (
            .O(N__28765),
            .I(N__28756));
    InMux I__6198 (
            .O(N__28764),
            .I(N__28756));
    InMux I__6197 (
            .O(N__28763),
            .I(N__28756));
    LocalMux I__6196 (
            .O(N__28756),
            .I(\this_ppu.N_329_0 ));
    CascadeMux I__6195 (
            .O(N__28753),
            .I(N__28750));
    CascadeBuf I__6194 (
            .O(N__28750),
            .I(N__28747));
    CascadeMux I__6193 (
            .O(N__28747),
            .I(N__28744));
    InMux I__6192 (
            .O(N__28744),
            .I(N__28741));
    LocalMux I__6191 (
            .O(N__28741),
            .I(N__28737));
    InMux I__6190 (
            .O(N__28740),
            .I(N__28730));
    Span4Mux_h I__6189 (
            .O(N__28737),
            .I(N__28724));
    InMux I__6188 (
            .O(N__28736),
            .I(N__28719));
    InMux I__6187 (
            .O(N__28735),
            .I(N__28719));
    InMux I__6186 (
            .O(N__28734),
            .I(N__28714));
    InMux I__6185 (
            .O(N__28733),
            .I(N__28714));
    LocalMux I__6184 (
            .O(N__28730),
            .I(N__28711));
    InMux I__6183 (
            .O(N__28729),
            .I(N__28706));
    InMux I__6182 (
            .O(N__28728),
            .I(N__28706));
    InMux I__6181 (
            .O(N__28727),
            .I(N__28703));
    Span4Mux_v I__6180 (
            .O(N__28724),
            .I(N__28700));
    LocalMux I__6179 (
            .O(N__28719),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__6178 (
            .O(N__28714),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__6177 (
            .O(N__28711),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__6176 (
            .O(N__28706),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__6175 (
            .O(N__28703),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__6174 (
            .O(N__28700),
            .I(M_this_ppu_oam_addr_0));
    CascadeMux I__6173 (
            .O(N__28687),
            .I(N__28684));
    CascadeBuf I__6172 (
            .O(N__28684),
            .I(N__28681));
    CascadeMux I__6171 (
            .O(N__28681),
            .I(N__28678));
    InMux I__6170 (
            .O(N__28678),
            .I(N__28675));
    LocalMux I__6169 (
            .O(N__28675),
            .I(N__28669));
    CascadeMux I__6168 (
            .O(N__28674),
            .I(N__28666));
    CascadeMux I__6167 (
            .O(N__28673),
            .I(N__28663));
    InMux I__6166 (
            .O(N__28672),
            .I(N__28658));
    Span4Mux_v I__6165 (
            .O(N__28669),
            .I(N__28654));
    InMux I__6164 (
            .O(N__28666),
            .I(N__28651));
    InMux I__6163 (
            .O(N__28663),
            .I(N__28648));
    InMux I__6162 (
            .O(N__28662),
            .I(N__28643));
    InMux I__6161 (
            .O(N__28661),
            .I(N__28643));
    LocalMux I__6160 (
            .O(N__28658),
            .I(N__28640));
    InMux I__6159 (
            .O(N__28657),
            .I(N__28637));
    Span4Mux_h I__6158 (
            .O(N__28654),
            .I(N__28634));
    LocalMux I__6157 (
            .O(N__28651),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__6156 (
            .O(N__28648),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__6155 (
            .O(N__28643),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__6154 (
            .O(N__28640),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__6153 (
            .O(N__28637),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__6152 (
            .O(N__28634),
            .I(M_this_ppu_oam_addr_1));
    InMux I__6151 (
            .O(N__28621),
            .I(N__28612));
    InMux I__6150 (
            .O(N__28620),
            .I(N__28612));
    InMux I__6149 (
            .O(N__28619),
            .I(N__28607));
    InMux I__6148 (
            .O(N__28618),
            .I(N__28607));
    InMux I__6147 (
            .O(N__28617),
            .I(N__28604));
    LocalMux I__6146 (
            .O(N__28612),
            .I(\this_ppu.un1_M_state_q_2_0 ));
    LocalMux I__6145 (
            .O(N__28607),
            .I(\this_ppu.un1_M_state_q_2_0 ));
    LocalMux I__6144 (
            .O(N__28604),
            .I(\this_ppu.un1_M_state_q_2_0 ));
    CascadeMux I__6143 (
            .O(N__28597),
            .I(N__28594));
    CascadeBuf I__6142 (
            .O(N__28594),
            .I(N__28591));
    CascadeMux I__6141 (
            .O(N__28591),
            .I(N__28588));
    InMux I__6140 (
            .O(N__28588),
            .I(N__28585));
    LocalMux I__6139 (
            .O(N__28585),
            .I(N__28582));
    Odrv12 I__6138 (
            .O(N__28582),
            .I(\this_ppu.N_19_0 ));
    CascadeMux I__6137 (
            .O(N__28579),
            .I(\this_ppu.un1_M_vaddress_q_c2_cascade_ ));
    InMux I__6136 (
            .O(N__28576),
            .I(N__28573));
    LocalMux I__6135 (
            .O(N__28573),
            .I(M_this_data_tmp_qZ0Z_8));
    InMux I__6134 (
            .O(N__28570),
            .I(N__28567));
    LocalMux I__6133 (
            .O(N__28567),
            .I(N__28564));
    Span4Mux_h I__6132 (
            .O(N__28564),
            .I(N__28561));
    Span4Mux_h I__6131 (
            .O(N__28561),
            .I(N__28558));
    Odrv4 I__6130 (
            .O(N__28558),
            .I(M_this_oam_ram_write_data_8));
    CascadeMux I__6129 (
            .O(N__28555),
            .I(\this_ppu.N_61_i_cascade_ ));
    CascadeMux I__6128 (
            .O(N__28552),
            .I(N__28549));
    InMux I__6127 (
            .O(N__28549),
            .I(N__28546));
    LocalMux I__6126 (
            .O(N__28546),
            .I(N__28542));
    InMux I__6125 (
            .O(N__28545),
            .I(N__28539));
    Span12Mux_h I__6124 (
            .O(N__28542),
            .I(N__28536));
    LocalMux I__6123 (
            .O(N__28539),
            .I(N__28533));
    Odrv12 I__6122 (
            .O(N__28536),
            .I(\this_ppu.N_769_0 ));
    Odrv4 I__6121 (
            .O(N__28533),
            .I(\this_ppu.N_769_0 ));
    InMux I__6120 (
            .O(N__28528),
            .I(N__28525));
    LocalMux I__6119 (
            .O(N__28525),
            .I(N__28522));
    Odrv4 I__6118 (
            .O(N__28522),
            .I(\this_ppu.M_state_q_srsts_i_i_o2_4_2 ));
    CascadeMux I__6117 (
            .O(N__28519),
            .I(N__28516));
    InMux I__6116 (
            .O(N__28516),
            .I(N__28512));
    InMux I__6115 (
            .O(N__28515),
            .I(N__28508));
    LocalMux I__6114 (
            .O(N__28512),
            .I(N__28504));
    InMux I__6113 (
            .O(N__28511),
            .I(N__28501));
    LocalMux I__6112 (
            .O(N__28508),
            .I(N__28498));
    InMux I__6111 (
            .O(N__28507),
            .I(N__28495));
    Span4Mux_h I__6110 (
            .O(N__28504),
            .I(N__28492));
    LocalMux I__6109 (
            .O(N__28501),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__6108 (
            .O(N__28498),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    LocalMux I__6107 (
            .O(N__28495),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__6106 (
            .O(N__28492),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    CascadeMux I__6105 (
            .O(N__28483),
            .I(\this_ppu.un1_M_state_q_2_0_cascade_ ));
    CascadeMux I__6104 (
            .O(N__28480),
            .I(N__28477));
    CascadeBuf I__6103 (
            .O(N__28477),
            .I(N__28474));
    CascadeMux I__6102 (
            .O(N__28474),
            .I(N__28471));
    InMux I__6101 (
            .O(N__28471),
            .I(N__28468));
    LocalMux I__6100 (
            .O(N__28468),
            .I(N__28465));
    Span4Mux_v I__6099 (
            .O(N__28465),
            .I(N__28459));
    InMux I__6098 (
            .O(N__28464),
            .I(N__28456));
    InMux I__6097 (
            .O(N__28463),
            .I(N__28453));
    InMux I__6096 (
            .O(N__28462),
            .I(N__28450));
    Span4Mux_h I__6095 (
            .O(N__28459),
            .I(N__28447));
    LocalMux I__6094 (
            .O(N__28456),
            .I(M_this_ppu_oam_addr_5));
    LocalMux I__6093 (
            .O(N__28453),
            .I(M_this_ppu_oam_addr_5));
    LocalMux I__6092 (
            .O(N__28450),
            .I(M_this_ppu_oam_addr_5));
    Odrv4 I__6091 (
            .O(N__28447),
            .I(M_this_ppu_oam_addr_5));
    InMux I__6090 (
            .O(N__28438),
            .I(N__28429));
    InMux I__6089 (
            .O(N__28437),
            .I(N__28426));
    InMux I__6088 (
            .O(N__28436),
            .I(N__28415));
    InMux I__6087 (
            .O(N__28435),
            .I(N__28415));
    InMux I__6086 (
            .O(N__28434),
            .I(N__28415));
    InMux I__6085 (
            .O(N__28433),
            .I(N__28415));
    InMux I__6084 (
            .O(N__28432),
            .I(N__28415));
    LocalMux I__6083 (
            .O(N__28429),
            .I(\this_ppu.M_oamcurr_qc_0_1 ));
    LocalMux I__6082 (
            .O(N__28426),
            .I(\this_ppu.M_oamcurr_qc_0_1 ));
    LocalMux I__6081 (
            .O(N__28415),
            .I(\this_ppu.M_oamcurr_qc_0_1 ));
    InMux I__6080 (
            .O(N__28408),
            .I(N__28404));
    InMux I__6079 (
            .O(N__28407),
            .I(N__28401));
    LocalMux I__6078 (
            .O(N__28404),
            .I(\this_ppu.un1_M_oamcurr_q_2_c5 ));
    LocalMux I__6077 (
            .O(N__28401),
            .I(\this_ppu.un1_M_oamcurr_q_2_c5 ));
    CascadeMux I__6076 (
            .O(N__28396),
            .I(N__28392));
    CascadeMux I__6075 (
            .O(N__28395),
            .I(N__28389));
    InMux I__6074 (
            .O(N__28392),
            .I(N__28384));
    InMux I__6073 (
            .O(N__28389),
            .I(N__28384));
    LocalMux I__6072 (
            .O(N__28384),
            .I(\this_ppu.M_oamcurr_qZ0Z_6 ));
    CascadeMux I__6071 (
            .O(N__28381),
            .I(N__28376));
    InMux I__6070 (
            .O(N__28380),
            .I(N__28372));
    InMux I__6069 (
            .O(N__28379),
            .I(N__28369));
    InMux I__6068 (
            .O(N__28376),
            .I(N__28366));
    InMux I__6067 (
            .O(N__28375),
            .I(N__28363));
    LocalMux I__6066 (
            .O(N__28372),
            .I(N__28360));
    LocalMux I__6065 (
            .O(N__28369),
            .I(N__28357));
    LocalMux I__6064 (
            .O(N__28366),
            .I(N__28353));
    LocalMux I__6063 (
            .O(N__28363),
            .I(N__28348));
    Span4Mux_v I__6062 (
            .O(N__28360),
            .I(N__28348));
    Span4Mux_v I__6061 (
            .O(N__28357),
            .I(N__28344));
    CascadeMux I__6060 (
            .O(N__28356),
            .I(N__28341));
    Span12Mux_s10_v I__6059 (
            .O(N__28353),
            .I(N__28338));
    Sp12to4 I__6058 (
            .O(N__28348),
            .I(N__28335));
    InMux I__6057 (
            .O(N__28347),
            .I(N__28332));
    Span4Mux_h I__6056 (
            .O(N__28344),
            .I(N__28329));
    InMux I__6055 (
            .O(N__28341),
            .I(N__28326));
    Odrv12 I__6054 (
            .O(N__28338),
            .I(M_this_ppu_vram_addr_2));
    Odrv12 I__6053 (
            .O(N__28335),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__6052 (
            .O(N__28332),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__6051 (
            .O(N__28329),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__6050 (
            .O(N__28326),
            .I(M_this_ppu_vram_addr_2));
    CascadeMux I__6049 (
            .O(N__28315),
            .I(N__28312));
    InMux I__6048 (
            .O(N__28312),
            .I(N__28309));
    LocalMux I__6047 (
            .O(N__28309),
            .I(M_this_scroll_qZ0Z_10));
    InMux I__6046 (
            .O(N__28306),
            .I(\this_ppu.un1_M_hoffset_d_cry_1 ));
    CascadeMux I__6045 (
            .O(N__28303),
            .I(N__28300));
    InMux I__6044 (
            .O(N__28300),
            .I(N__28296));
    InMux I__6043 (
            .O(N__28299),
            .I(N__28292));
    LocalMux I__6042 (
            .O(N__28296),
            .I(N__28289));
    CascadeMux I__6041 (
            .O(N__28295),
            .I(N__28286));
    LocalMux I__6040 (
            .O(N__28292),
            .I(N__28282));
    Span4Mux_h I__6039 (
            .O(N__28289),
            .I(N__28279));
    InMux I__6038 (
            .O(N__28286),
            .I(N__28272));
    InMux I__6037 (
            .O(N__28285),
            .I(N__28269));
    Span4Mux_v I__6036 (
            .O(N__28282),
            .I(N__28266));
    Span4Mux_h I__6035 (
            .O(N__28279),
            .I(N__28263));
    InMux I__6034 (
            .O(N__28278),
            .I(N__28260));
    InMux I__6033 (
            .O(N__28277),
            .I(N__28257));
    InMux I__6032 (
            .O(N__28276),
            .I(N__28254));
    InMux I__6031 (
            .O(N__28275),
            .I(N__28251));
    LocalMux I__6030 (
            .O(N__28272),
            .I(N__28246));
    LocalMux I__6029 (
            .O(N__28269),
            .I(N__28246));
    Span4Mux_h I__6028 (
            .O(N__28266),
            .I(N__28243));
    Span4Mux_v I__6027 (
            .O(N__28263),
            .I(N__28236));
    LocalMux I__6026 (
            .O(N__28260),
            .I(N__28236));
    LocalMux I__6025 (
            .O(N__28257),
            .I(N__28236));
    LocalMux I__6024 (
            .O(N__28254),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__6023 (
            .O(N__28251),
            .I(M_this_ppu_vram_addr_3));
    Odrv4 I__6022 (
            .O(N__28246),
            .I(M_this_ppu_vram_addr_3));
    Odrv4 I__6021 (
            .O(N__28243),
            .I(M_this_ppu_vram_addr_3));
    Odrv4 I__6020 (
            .O(N__28236),
            .I(M_this_ppu_vram_addr_3));
    CascadeMux I__6019 (
            .O(N__28225),
            .I(N__28222));
    InMux I__6018 (
            .O(N__28222),
            .I(N__28219));
    LocalMux I__6017 (
            .O(N__28219),
            .I(M_this_scroll_qZ0Z_11));
    InMux I__6016 (
            .O(N__28216),
            .I(\this_ppu.un1_M_hoffset_d_cry_2 ));
    CascadeMux I__6015 (
            .O(N__28213),
            .I(N__28210));
    InMux I__6014 (
            .O(N__28210),
            .I(N__28207));
    LocalMux I__6013 (
            .O(N__28207),
            .I(N__28203));
    InMux I__6012 (
            .O(N__28206),
            .I(N__28200));
    Span4Mux_h I__6011 (
            .O(N__28203),
            .I(N__28197));
    LocalMux I__6010 (
            .O(N__28200),
            .I(N__28191));
    Span4Mux_v I__6009 (
            .O(N__28197),
            .I(N__28188));
    CascadeMux I__6008 (
            .O(N__28196),
            .I(N__28185));
    InMux I__6007 (
            .O(N__28195),
            .I(N__28180));
    InMux I__6006 (
            .O(N__28194),
            .I(N__28180));
    Span4Mux_v I__6005 (
            .O(N__28191),
            .I(N__28177));
    Span4Mux_h I__6004 (
            .O(N__28188),
            .I(N__28174));
    InMux I__6003 (
            .O(N__28185),
            .I(N__28171));
    LocalMux I__6002 (
            .O(N__28180),
            .I(N__28166));
    Span4Mux_h I__6001 (
            .O(N__28177),
            .I(N__28166));
    Odrv4 I__6000 (
            .O(N__28174),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__5999 (
            .O(N__28171),
            .I(M_this_ppu_vram_addr_4));
    Odrv4 I__5998 (
            .O(N__28166),
            .I(M_this_ppu_vram_addr_4));
    CascadeMux I__5997 (
            .O(N__28159),
            .I(N__28156));
    InMux I__5996 (
            .O(N__28156),
            .I(N__28153));
    LocalMux I__5995 (
            .O(N__28153),
            .I(N__28150));
    Odrv4 I__5994 (
            .O(N__28150),
            .I(M_this_scroll_qZ0Z_12));
    InMux I__5993 (
            .O(N__28147),
            .I(\this_ppu.un1_M_hoffset_d_cry_3 ));
    InMux I__5992 (
            .O(N__28144),
            .I(N__28141));
    LocalMux I__5991 (
            .O(N__28141),
            .I(M_this_scroll_qZ0Z_13));
    CascadeMux I__5990 (
            .O(N__28138),
            .I(N__28135));
    InMux I__5989 (
            .O(N__28135),
            .I(N__28132));
    LocalMux I__5988 (
            .O(N__28132),
            .I(N__28128));
    CascadeMux I__5987 (
            .O(N__28131),
            .I(N__28125));
    Span4Mux_h I__5986 (
            .O(N__28128),
            .I(N__28122));
    InMux I__5985 (
            .O(N__28125),
            .I(N__28119));
    Span4Mux_h I__5984 (
            .O(N__28122),
            .I(N__28114));
    LocalMux I__5983 (
            .O(N__28119),
            .I(N__28111));
    InMux I__5982 (
            .O(N__28118),
            .I(N__28106));
    InMux I__5981 (
            .O(N__28117),
            .I(N__28106));
    Sp12to4 I__5980 (
            .O(N__28114),
            .I(N__28101));
    Span12Mux_h I__5979 (
            .O(N__28111),
            .I(N__28101));
    LocalMux I__5978 (
            .O(N__28106),
            .I(M_this_ppu_vram_addr_5));
    Odrv12 I__5977 (
            .O(N__28101),
            .I(M_this_ppu_vram_addr_5));
    InMux I__5976 (
            .O(N__28096),
            .I(\this_ppu.un1_M_hoffset_d_cry_4 ));
    InMux I__5975 (
            .O(N__28093),
            .I(N__28090));
    LocalMux I__5974 (
            .O(N__28090),
            .I(M_this_scroll_qZ0Z_14));
    CascadeMux I__5973 (
            .O(N__28087),
            .I(N__28083));
    CascadeMux I__5972 (
            .O(N__28086),
            .I(N__28080));
    InMux I__5971 (
            .O(N__28083),
            .I(N__28077));
    InMux I__5970 (
            .O(N__28080),
            .I(N__28074));
    LocalMux I__5969 (
            .O(N__28077),
            .I(N__28071));
    LocalMux I__5968 (
            .O(N__28074),
            .I(N__28068));
    Sp12to4 I__5967 (
            .O(N__28071),
            .I(N__28063));
    Span4Mux_v I__5966 (
            .O(N__28068),
            .I(N__28060));
    InMux I__5965 (
            .O(N__28067),
            .I(N__28057));
    InMux I__5964 (
            .O(N__28066),
            .I(N__28054));
    Span12Mux_s9_v I__5963 (
            .O(N__28063),
            .I(N__28051));
    Span4Mux_h I__5962 (
            .O(N__28060),
            .I(N__28048));
    LocalMux I__5961 (
            .O(N__28057),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__5960 (
            .O(N__28054),
            .I(M_this_ppu_vram_addr_6));
    Odrv12 I__5959 (
            .O(N__28051),
            .I(M_this_ppu_vram_addr_6));
    Odrv4 I__5958 (
            .O(N__28048),
            .I(M_this_ppu_vram_addr_6));
    InMux I__5957 (
            .O(N__28039),
            .I(\this_ppu.un1_M_hoffset_d_cry_5 ));
    InMux I__5956 (
            .O(N__28036),
            .I(N__28033));
    LocalMux I__5955 (
            .O(N__28033),
            .I(N__28029));
    InMux I__5954 (
            .O(N__28032),
            .I(N__28026));
    Span4Mux_v I__5953 (
            .O(N__28029),
            .I(N__28023));
    LocalMux I__5952 (
            .O(N__28026),
            .I(N__28018));
    Span4Mux_v I__5951 (
            .O(N__28023),
            .I(N__28018));
    Odrv4 I__5950 (
            .O(N__28018),
            .I(\this_ppu.M_haddress_qZ0Z_7 ));
    CascadeMux I__5949 (
            .O(N__28015),
            .I(N__28012));
    InMux I__5948 (
            .O(N__28012),
            .I(N__28009));
    LocalMux I__5947 (
            .O(N__28009),
            .I(M_this_scroll_qZ0Z_15));
    InMux I__5946 (
            .O(N__28006),
            .I(\this_ppu.un1_M_hoffset_d_cry_6 ));
    InMux I__5945 (
            .O(N__28003),
            .I(bfn_19_18_0_));
    InMux I__5944 (
            .O(N__28000),
            .I(N__27997));
    LocalMux I__5943 (
            .O(N__27997),
            .I(N__27994));
    Span4Mux_h I__5942 (
            .O(N__27994),
            .I(N__27991));
    Span4Mux_h I__5941 (
            .O(N__27991),
            .I(N__27988));
    Odrv4 I__5940 (
            .O(N__27988),
            .I(\this_ppu.oam_cache.mem_1 ));
    InMux I__5939 (
            .O(N__27985),
            .I(N__27982));
    LocalMux I__5938 (
            .O(N__27982),
            .I(N__27979));
    Span4Mux_h I__5937 (
            .O(N__27979),
            .I(N__27976));
    Odrv4 I__5936 (
            .O(N__27976),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_1 ));
    CEMux I__5935 (
            .O(N__27973),
            .I(N__27969));
    CEMux I__5934 (
            .O(N__27972),
            .I(N__27966));
    LocalMux I__5933 (
            .O(N__27969),
            .I(N_1310_0));
    LocalMux I__5932 (
            .O(N__27966),
            .I(N_1310_0));
    CascadeMux I__5931 (
            .O(N__27961),
            .I(N__27958));
    InMux I__5930 (
            .O(N__27958),
            .I(N__27955));
    LocalMux I__5929 (
            .O(N__27955),
            .I(N__27951));
    InMux I__5928 (
            .O(N__27954),
            .I(N__27948));
    Sp12to4 I__5927 (
            .O(N__27951),
            .I(N__27945));
    LocalMux I__5926 (
            .O(N__27948),
            .I(N__27939));
    Span12Mux_h I__5925 (
            .O(N__27945),
            .I(N__27935));
    InMux I__5924 (
            .O(N__27944),
            .I(N__27930));
    InMux I__5923 (
            .O(N__27943),
            .I(N__27930));
    InMux I__5922 (
            .O(N__27942),
            .I(N__27927));
    Span12Mux_v I__5921 (
            .O(N__27939),
            .I(N__27924));
    InMux I__5920 (
            .O(N__27938),
            .I(N__27921));
    Odrv12 I__5919 (
            .O(N__27935),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__5918 (
            .O(N__27930),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__5917 (
            .O(N__27927),
            .I(M_this_ppu_vram_addr_1));
    Odrv12 I__5916 (
            .O(N__27924),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__5915 (
            .O(N__27921),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__5914 (
            .O(N__27910),
            .I(N__27907));
    InMux I__5913 (
            .O(N__27907),
            .I(N__27904));
    LocalMux I__5912 (
            .O(N__27904),
            .I(M_this_scroll_qZ0Z_9));
    InMux I__5911 (
            .O(N__27901),
            .I(\this_ppu.un1_M_hoffset_d_cry_0 ));
    CascadeMux I__5910 (
            .O(N__27898),
            .I(N__27894));
    CascadeMux I__5909 (
            .O(N__27897),
            .I(N__27889));
    InMux I__5908 (
            .O(N__27894),
            .I(N__27884));
    CascadeMux I__5907 (
            .O(N__27893),
            .I(N__27881));
    CascadeMux I__5906 (
            .O(N__27892),
            .I(N__27876));
    InMux I__5905 (
            .O(N__27889),
            .I(N__27872));
    CascadeMux I__5904 (
            .O(N__27888),
            .I(N__27869));
    CascadeMux I__5903 (
            .O(N__27887),
            .I(N__27865));
    LocalMux I__5902 (
            .O(N__27884),
            .I(N__27862));
    InMux I__5901 (
            .O(N__27881),
            .I(N__27859));
    CascadeMux I__5900 (
            .O(N__27880),
            .I(N__27856));
    CascadeMux I__5899 (
            .O(N__27879),
            .I(N__27848));
    InMux I__5898 (
            .O(N__27876),
            .I(N__27844));
    CascadeMux I__5897 (
            .O(N__27875),
            .I(N__27841));
    LocalMux I__5896 (
            .O(N__27872),
            .I(N__27838));
    InMux I__5895 (
            .O(N__27869),
            .I(N__27835));
    CascadeMux I__5894 (
            .O(N__27868),
            .I(N__27832));
    InMux I__5893 (
            .O(N__27865),
            .I(N__27829));
    Span4Mux_h I__5892 (
            .O(N__27862),
            .I(N__27826));
    LocalMux I__5891 (
            .O(N__27859),
            .I(N__27823));
    InMux I__5890 (
            .O(N__27856),
            .I(N__27820));
    CascadeMux I__5889 (
            .O(N__27855),
            .I(N__27817));
    CascadeMux I__5888 (
            .O(N__27854),
            .I(N__27814));
    CascadeMux I__5887 (
            .O(N__27853),
            .I(N__27811));
    CascadeMux I__5886 (
            .O(N__27852),
            .I(N__27808));
    CascadeMux I__5885 (
            .O(N__27851),
            .I(N__27805));
    InMux I__5884 (
            .O(N__27848),
            .I(N__27802));
    CascadeMux I__5883 (
            .O(N__27847),
            .I(N__27799));
    LocalMux I__5882 (
            .O(N__27844),
            .I(N__27796));
    InMux I__5881 (
            .O(N__27841),
            .I(N__27793));
    Span4Mux_h I__5880 (
            .O(N__27838),
            .I(N__27790));
    LocalMux I__5879 (
            .O(N__27835),
            .I(N__27787));
    InMux I__5878 (
            .O(N__27832),
            .I(N__27784));
    LocalMux I__5877 (
            .O(N__27829),
            .I(N__27781));
    Span4Mux_v I__5876 (
            .O(N__27826),
            .I(N__27776));
    Span4Mux_h I__5875 (
            .O(N__27823),
            .I(N__27776));
    LocalMux I__5874 (
            .O(N__27820),
            .I(N__27773));
    InMux I__5873 (
            .O(N__27817),
            .I(N__27770));
    InMux I__5872 (
            .O(N__27814),
            .I(N__27767));
    InMux I__5871 (
            .O(N__27811),
            .I(N__27764));
    InMux I__5870 (
            .O(N__27808),
            .I(N__27761));
    InMux I__5869 (
            .O(N__27805),
            .I(N__27758));
    LocalMux I__5868 (
            .O(N__27802),
            .I(N__27755));
    InMux I__5867 (
            .O(N__27799),
            .I(N__27752));
    Span4Mux_h I__5866 (
            .O(N__27796),
            .I(N__27749));
    LocalMux I__5865 (
            .O(N__27793),
            .I(N__27746));
    Span4Mux_v I__5864 (
            .O(N__27790),
            .I(N__27741));
    Span4Mux_h I__5863 (
            .O(N__27787),
            .I(N__27741));
    LocalMux I__5862 (
            .O(N__27784),
            .I(N__27738));
    Span4Mux_h I__5861 (
            .O(N__27781),
            .I(N__27735));
    Span4Mux_v I__5860 (
            .O(N__27776),
            .I(N__27730));
    Span4Mux_h I__5859 (
            .O(N__27773),
            .I(N__27730));
    LocalMux I__5858 (
            .O(N__27770),
            .I(N__27727));
    LocalMux I__5857 (
            .O(N__27767),
            .I(N__27718));
    LocalMux I__5856 (
            .O(N__27764),
            .I(N__27718));
    LocalMux I__5855 (
            .O(N__27761),
            .I(N__27718));
    LocalMux I__5854 (
            .O(N__27758),
            .I(N__27718));
    Sp12to4 I__5853 (
            .O(N__27755),
            .I(N__27713));
    LocalMux I__5852 (
            .O(N__27752),
            .I(N__27713));
    Span4Mux_v I__5851 (
            .O(N__27749),
            .I(N__27708));
    Span4Mux_h I__5850 (
            .O(N__27746),
            .I(N__27708));
    Span4Mux_v I__5849 (
            .O(N__27741),
            .I(N__27703));
    Span4Mux_h I__5848 (
            .O(N__27738),
            .I(N__27703));
    Span4Mux_v I__5847 (
            .O(N__27735),
            .I(N__27696));
    Span4Mux_v I__5846 (
            .O(N__27730),
            .I(N__27696));
    Span4Mux_h I__5845 (
            .O(N__27727),
            .I(N__27696));
    Span12Mux_v I__5844 (
            .O(N__27718),
            .I(N__27690));
    Span12Mux_v I__5843 (
            .O(N__27713),
            .I(N__27690));
    Span4Mux_h I__5842 (
            .O(N__27708),
            .I(N__27685));
    Span4Mux_h I__5841 (
            .O(N__27703),
            .I(N__27685));
    Span4Mux_h I__5840 (
            .O(N__27696),
            .I(N__27682));
    InMux I__5839 (
            .O(N__27695),
            .I(N__27679));
    Odrv12 I__5838 (
            .O(N__27690),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv4 I__5837 (
            .O(N__27685),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv4 I__5836 (
            .O(N__27682),
            .I(M_this_spr_address_qZ0Z_7));
    LocalMux I__5835 (
            .O(N__27679),
            .I(M_this_spr_address_qZ0Z_7));
    InMux I__5834 (
            .O(N__27670),
            .I(un1_M_this_spr_address_q_cry_6));
    CascadeMux I__5833 (
            .O(N__27667),
            .I(N__27663));
    CascadeMux I__5832 (
            .O(N__27666),
            .I(N__27659));
    InMux I__5831 (
            .O(N__27663),
            .I(N__27655));
    CascadeMux I__5830 (
            .O(N__27662),
            .I(N__27652));
    InMux I__5829 (
            .O(N__27659),
            .I(N__27647));
    CascadeMux I__5828 (
            .O(N__27658),
            .I(N__27644));
    LocalMux I__5827 (
            .O(N__27655),
            .I(N__27639));
    InMux I__5826 (
            .O(N__27652),
            .I(N__27636));
    CascadeMux I__5825 (
            .O(N__27651),
            .I(N__27633));
    CascadeMux I__5824 (
            .O(N__27650),
            .I(N__27630));
    LocalMux I__5823 (
            .O(N__27647),
            .I(N__27626));
    InMux I__5822 (
            .O(N__27644),
            .I(N__27623));
    CascadeMux I__5821 (
            .O(N__27643),
            .I(N__27620));
    CascadeMux I__5820 (
            .O(N__27642),
            .I(N__27616));
    Span4Mux_h I__5819 (
            .O(N__27639),
            .I(N__27606));
    LocalMux I__5818 (
            .O(N__27636),
            .I(N__27606));
    InMux I__5817 (
            .O(N__27633),
            .I(N__27603));
    InMux I__5816 (
            .O(N__27630),
            .I(N__27600));
    CascadeMux I__5815 (
            .O(N__27629),
            .I(N__27597));
    Span4Mux_v I__5814 (
            .O(N__27626),
            .I(N__27592));
    LocalMux I__5813 (
            .O(N__27623),
            .I(N__27592));
    InMux I__5812 (
            .O(N__27620),
            .I(N__27589));
    CascadeMux I__5811 (
            .O(N__27619),
            .I(N__27586));
    InMux I__5810 (
            .O(N__27616),
            .I(N__27583));
    CascadeMux I__5809 (
            .O(N__27615),
            .I(N__27580));
    CascadeMux I__5808 (
            .O(N__27614),
            .I(N__27577));
    CascadeMux I__5807 (
            .O(N__27613),
            .I(N__27574));
    CascadeMux I__5806 (
            .O(N__27612),
            .I(N__27571));
    CascadeMux I__5805 (
            .O(N__27611),
            .I(N__27568));
    Span4Mux_v I__5804 (
            .O(N__27606),
            .I(N__27563));
    LocalMux I__5803 (
            .O(N__27603),
            .I(N__27563));
    LocalMux I__5802 (
            .O(N__27600),
            .I(N__27560));
    InMux I__5801 (
            .O(N__27597),
            .I(N__27557));
    Span4Mux_h I__5800 (
            .O(N__27592),
            .I(N__27552));
    LocalMux I__5799 (
            .O(N__27589),
            .I(N__27552));
    InMux I__5798 (
            .O(N__27586),
            .I(N__27549));
    LocalMux I__5797 (
            .O(N__27583),
            .I(N__27546));
    InMux I__5796 (
            .O(N__27580),
            .I(N__27543));
    InMux I__5795 (
            .O(N__27577),
            .I(N__27540));
    InMux I__5794 (
            .O(N__27574),
            .I(N__27536));
    InMux I__5793 (
            .O(N__27571),
            .I(N__27533));
    InMux I__5792 (
            .O(N__27568),
            .I(N__27530));
    Span4Mux_v I__5791 (
            .O(N__27563),
            .I(N__27525));
    Span4Mux_v I__5790 (
            .O(N__27560),
            .I(N__27525));
    LocalMux I__5789 (
            .O(N__27557),
            .I(N__27522));
    Span4Mux_v I__5788 (
            .O(N__27552),
            .I(N__27517));
    LocalMux I__5787 (
            .O(N__27549),
            .I(N__27517));
    Span4Mux_v I__5786 (
            .O(N__27546),
            .I(N__27510));
    LocalMux I__5785 (
            .O(N__27543),
            .I(N__27510));
    LocalMux I__5784 (
            .O(N__27540),
            .I(N__27510));
    CascadeMux I__5783 (
            .O(N__27539),
            .I(N__27507));
    LocalMux I__5782 (
            .O(N__27536),
            .I(N__27504));
    LocalMux I__5781 (
            .O(N__27533),
            .I(N__27501));
    LocalMux I__5780 (
            .O(N__27530),
            .I(N__27498));
    Sp12to4 I__5779 (
            .O(N__27525),
            .I(N__27493));
    Sp12to4 I__5778 (
            .O(N__27522),
            .I(N__27493));
    Span4Mux_v I__5777 (
            .O(N__27517),
            .I(N__27488));
    Span4Mux_v I__5776 (
            .O(N__27510),
            .I(N__27488));
    InMux I__5775 (
            .O(N__27507),
            .I(N__27485));
    Span12Mux_h I__5774 (
            .O(N__27504),
            .I(N__27481));
    Span12Mux_h I__5773 (
            .O(N__27501),
            .I(N__27476));
    Span12Mux_h I__5772 (
            .O(N__27498),
            .I(N__27476));
    Span12Mux_h I__5771 (
            .O(N__27493),
            .I(N__27469));
    Sp12to4 I__5770 (
            .O(N__27488),
            .I(N__27469));
    LocalMux I__5769 (
            .O(N__27485),
            .I(N__27469));
    InMux I__5768 (
            .O(N__27484),
            .I(N__27466));
    Odrv12 I__5767 (
            .O(N__27481),
            .I(M_this_spr_address_qZ0Z_8));
    Odrv12 I__5766 (
            .O(N__27476),
            .I(M_this_spr_address_qZ0Z_8));
    Odrv12 I__5765 (
            .O(N__27469),
            .I(M_this_spr_address_qZ0Z_8));
    LocalMux I__5764 (
            .O(N__27466),
            .I(M_this_spr_address_qZ0Z_8));
    InMux I__5763 (
            .O(N__27457),
            .I(bfn_19_14_0_));
    CascadeMux I__5762 (
            .O(N__27454),
            .I(N__27450));
    CascadeMux I__5761 (
            .O(N__27453),
            .I(N__27446));
    InMux I__5760 (
            .O(N__27450),
            .I(N__27442));
    CascadeMux I__5759 (
            .O(N__27449),
            .I(N__27439));
    InMux I__5758 (
            .O(N__27446),
            .I(N__27435));
    CascadeMux I__5757 (
            .O(N__27445),
            .I(N__27432));
    LocalMux I__5756 (
            .O(N__27442),
            .I(N__27428));
    InMux I__5755 (
            .O(N__27439),
            .I(N__27425));
    CascadeMux I__5754 (
            .O(N__27438),
            .I(N__27422));
    LocalMux I__5753 (
            .O(N__27435),
            .I(N__27417));
    InMux I__5752 (
            .O(N__27432),
            .I(N__27414));
    CascadeMux I__5751 (
            .O(N__27431),
            .I(N__27411));
    Span4Mux_h I__5750 (
            .O(N__27428),
            .I(N__27403));
    LocalMux I__5749 (
            .O(N__27425),
            .I(N__27403));
    InMux I__5748 (
            .O(N__27422),
            .I(N__27400));
    CascadeMux I__5747 (
            .O(N__27421),
            .I(N__27397));
    CascadeMux I__5746 (
            .O(N__27420),
            .I(N__27394));
    Span4Mux_v I__5745 (
            .O(N__27417),
            .I(N__27388));
    LocalMux I__5744 (
            .O(N__27414),
            .I(N__27388));
    InMux I__5743 (
            .O(N__27411),
            .I(N__27385));
    CascadeMux I__5742 (
            .O(N__27410),
            .I(N__27382));
    CascadeMux I__5741 (
            .O(N__27409),
            .I(N__27378));
    CascadeMux I__5740 (
            .O(N__27408),
            .I(N__27373));
    Span4Mux_v I__5739 (
            .O(N__27403),
            .I(N__27368));
    LocalMux I__5738 (
            .O(N__27400),
            .I(N__27368));
    InMux I__5737 (
            .O(N__27397),
            .I(N__27365));
    InMux I__5736 (
            .O(N__27394),
            .I(N__27362));
    CascadeMux I__5735 (
            .O(N__27393),
            .I(N__27359));
    Span4Mux_h I__5734 (
            .O(N__27388),
            .I(N__27354));
    LocalMux I__5733 (
            .O(N__27385),
            .I(N__27354));
    InMux I__5732 (
            .O(N__27382),
            .I(N__27351));
    CascadeMux I__5731 (
            .O(N__27381),
            .I(N__27348));
    InMux I__5730 (
            .O(N__27378),
            .I(N__27345));
    CascadeMux I__5729 (
            .O(N__27377),
            .I(N__27342));
    CascadeMux I__5728 (
            .O(N__27376),
            .I(N__27339));
    InMux I__5727 (
            .O(N__27373),
            .I(N__27336));
    Span4Mux_h I__5726 (
            .O(N__27368),
            .I(N__27331));
    LocalMux I__5725 (
            .O(N__27365),
            .I(N__27331));
    LocalMux I__5724 (
            .O(N__27362),
            .I(N__27328));
    InMux I__5723 (
            .O(N__27359),
            .I(N__27325));
    Span4Mux_v I__5722 (
            .O(N__27354),
            .I(N__27320));
    LocalMux I__5721 (
            .O(N__27351),
            .I(N__27320));
    InMux I__5720 (
            .O(N__27348),
            .I(N__27317));
    LocalMux I__5719 (
            .O(N__27345),
            .I(N__27314));
    InMux I__5718 (
            .O(N__27342),
            .I(N__27311));
    InMux I__5717 (
            .O(N__27339),
            .I(N__27308));
    LocalMux I__5716 (
            .O(N__27336),
            .I(N__27304));
    Span4Mux_v I__5715 (
            .O(N__27331),
            .I(N__27297));
    Span4Mux_v I__5714 (
            .O(N__27328),
            .I(N__27297));
    LocalMux I__5713 (
            .O(N__27325),
            .I(N__27297));
    Span4Mux_h I__5712 (
            .O(N__27320),
            .I(N__27292));
    LocalMux I__5711 (
            .O(N__27317),
            .I(N__27292));
    Span4Mux_v I__5710 (
            .O(N__27314),
            .I(N__27285));
    LocalMux I__5709 (
            .O(N__27311),
            .I(N__27285));
    LocalMux I__5708 (
            .O(N__27308),
            .I(N__27285));
    CascadeMux I__5707 (
            .O(N__27307),
            .I(N__27282));
    Span12Mux_h I__5706 (
            .O(N__27304),
            .I(N__27279));
    Sp12to4 I__5705 (
            .O(N__27297),
            .I(N__27276));
    Span4Mux_v I__5704 (
            .O(N__27292),
            .I(N__27271));
    Span4Mux_v I__5703 (
            .O(N__27285),
            .I(N__27271));
    InMux I__5702 (
            .O(N__27282),
            .I(N__27268));
    Span12Mux_v I__5701 (
            .O(N__27279),
            .I(N__27258));
    Span12Mux_h I__5700 (
            .O(N__27276),
            .I(N__27258));
    Sp12to4 I__5699 (
            .O(N__27271),
            .I(N__27258));
    LocalMux I__5698 (
            .O(N__27268),
            .I(N__27258));
    InMux I__5697 (
            .O(N__27267),
            .I(N__27255));
    Odrv12 I__5696 (
            .O(N__27258),
            .I(M_this_spr_address_qZ0Z_9));
    LocalMux I__5695 (
            .O(N__27255),
            .I(M_this_spr_address_qZ0Z_9));
    InMux I__5694 (
            .O(N__27250),
            .I(un1_M_this_spr_address_q_cry_8));
    CascadeMux I__5693 (
            .O(N__27247),
            .I(N__27244));
    InMux I__5692 (
            .O(N__27244),
            .I(N__27240));
    CascadeMux I__5691 (
            .O(N__27243),
            .I(N__27237));
    LocalMux I__5690 (
            .O(N__27240),
            .I(N__27230));
    InMux I__5689 (
            .O(N__27237),
            .I(N__27227));
    CascadeMux I__5688 (
            .O(N__27236),
            .I(N__27224));
    CascadeMux I__5687 (
            .O(N__27235),
            .I(N__27218));
    CascadeMux I__5686 (
            .O(N__27234),
            .I(N__27215));
    CascadeMux I__5685 (
            .O(N__27233),
            .I(N__27210));
    Span4Mux_h I__5684 (
            .O(N__27230),
            .I(N__27204));
    LocalMux I__5683 (
            .O(N__27227),
            .I(N__27204));
    InMux I__5682 (
            .O(N__27224),
            .I(N__27201));
    CascadeMux I__5681 (
            .O(N__27223),
            .I(N__27198));
    CascadeMux I__5680 (
            .O(N__27222),
            .I(N__27195));
    CascadeMux I__5679 (
            .O(N__27221),
            .I(N__27190));
    InMux I__5678 (
            .O(N__27218),
            .I(N__27187));
    InMux I__5677 (
            .O(N__27215),
            .I(N__27183));
    CascadeMux I__5676 (
            .O(N__27214),
            .I(N__27180));
    CascadeMux I__5675 (
            .O(N__27213),
            .I(N__27177));
    InMux I__5674 (
            .O(N__27210),
            .I(N__27173));
    CascadeMux I__5673 (
            .O(N__27209),
            .I(N__27170));
    Span4Mux_v I__5672 (
            .O(N__27204),
            .I(N__27165));
    LocalMux I__5671 (
            .O(N__27201),
            .I(N__27165));
    InMux I__5670 (
            .O(N__27198),
            .I(N__27162));
    InMux I__5669 (
            .O(N__27195),
            .I(N__27159));
    CascadeMux I__5668 (
            .O(N__27194),
            .I(N__27156));
    CascadeMux I__5667 (
            .O(N__27193),
            .I(N__27153));
    InMux I__5666 (
            .O(N__27190),
            .I(N__27150));
    LocalMux I__5665 (
            .O(N__27187),
            .I(N__27147));
    CascadeMux I__5664 (
            .O(N__27186),
            .I(N__27144));
    LocalMux I__5663 (
            .O(N__27183),
            .I(N__27141));
    InMux I__5662 (
            .O(N__27180),
            .I(N__27138));
    InMux I__5661 (
            .O(N__27177),
            .I(N__27135));
    CascadeMux I__5660 (
            .O(N__27176),
            .I(N__27132));
    LocalMux I__5659 (
            .O(N__27173),
            .I(N__27129));
    InMux I__5658 (
            .O(N__27170),
            .I(N__27126));
    Span4Mux_h I__5657 (
            .O(N__27165),
            .I(N__27123));
    LocalMux I__5656 (
            .O(N__27162),
            .I(N__27120));
    LocalMux I__5655 (
            .O(N__27159),
            .I(N__27117));
    InMux I__5654 (
            .O(N__27156),
            .I(N__27114));
    InMux I__5653 (
            .O(N__27153),
            .I(N__27111));
    LocalMux I__5652 (
            .O(N__27150),
            .I(N__27108));
    Span4Mux_v I__5651 (
            .O(N__27147),
            .I(N__27105));
    InMux I__5650 (
            .O(N__27144),
            .I(N__27102));
    Span4Mux_h I__5649 (
            .O(N__27141),
            .I(N__27099));
    LocalMux I__5648 (
            .O(N__27138),
            .I(N__27096));
    LocalMux I__5647 (
            .O(N__27135),
            .I(N__27093));
    InMux I__5646 (
            .O(N__27132),
            .I(N__27090));
    Span12Mux_s1_v I__5645 (
            .O(N__27129),
            .I(N__27085));
    LocalMux I__5644 (
            .O(N__27126),
            .I(N__27085));
    Span4Mux_v I__5643 (
            .O(N__27123),
            .I(N__27080));
    Span4Mux_h I__5642 (
            .O(N__27120),
            .I(N__27080));
    Sp12to4 I__5641 (
            .O(N__27117),
            .I(N__27077));
    LocalMux I__5640 (
            .O(N__27114),
            .I(N__27074));
    LocalMux I__5639 (
            .O(N__27111),
            .I(N__27071));
    Span12Mux_h I__5638 (
            .O(N__27108),
            .I(N__27064));
    Sp12to4 I__5637 (
            .O(N__27105),
            .I(N__27064));
    LocalMux I__5636 (
            .O(N__27102),
            .I(N__27064));
    Span4Mux_v I__5635 (
            .O(N__27099),
            .I(N__27059));
    Span4Mux_h I__5634 (
            .O(N__27096),
            .I(N__27059));
    Span4Mux_h I__5633 (
            .O(N__27093),
            .I(N__27056));
    LocalMux I__5632 (
            .O(N__27090),
            .I(N__27053));
    Span12Mux_v I__5631 (
            .O(N__27085),
            .I(N__27049));
    Span4Mux_h I__5630 (
            .O(N__27080),
            .I(N__27046));
    Span12Mux_h I__5629 (
            .O(N__27077),
            .I(N__27041));
    Span12Mux_h I__5628 (
            .O(N__27074),
            .I(N__27041));
    Span12Mux_h I__5627 (
            .O(N__27071),
            .I(N__27036));
    Span12Mux_h I__5626 (
            .O(N__27064),
            .I(N__27036));
    Span4Mux_v I__5625 (
            .O(N__27059),
            .I(N__27029));
    Span4Mux_v I__5624 (
            .O(N__27056),
            .I(N__27029));
    Span4Mux_h I__5623 (
            .O(N__27053),
            .I(N__27029));
    InMux I__5622 (
            .O(N__27052),
            .I(N__27026));
    Odrv12 I__5621 (
            .O(N__27049),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv4 I__5620 (
            .O(N__27046),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv12 I__5619 (
            .O(N__27041),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv12 I__5618 (
            .O(N__27036),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv4 I__5617 (
            .O(N__27029),
            .I(M_this_spr_address_qZ0Z_10));
    LocalMux I__5616 (
            .O(N__27026),
            .I(M_this_spr_address_qZ0Z_10));
    InMux I__5615 (
            .O(N__27013),
            .I(un1_M_this_spr_address_q_cry_9));
    InMux I__5614 (
            .O(N__27010),
            .I(un1_M_this_spr_address_q_cry_10));
    InMux I__5613 (
            .O(N__27007),
            .I(un1_M_this_spr_address_q_cry_11));
    InMux I__5612 (
            .O(N__27004),
            .I(un1_M_this_spr_address_q_cry_12));
    InMux I__5611 (
            .O(N__27001),
            .I(N__26998));
    LocalMux I__5610 (
            .O(N__26998),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__5609 (
            .O(N__26995),
            .I(N__26992));
    LocalMux I__5608 (
            .O(N__26992),
            .I(N__26989));
    Span4Mux_h I__5607 (
            .O(N__26989),
            .I(N__26986));
    Span4Mux_h I__5606 (
            .O(N__26986),
            .I(N__26983));
    Odrv4 I__5605 (
            .O(N__26983),
            .I(M_this_oam_ram_write_data_18));
    InMux I__5604 (
            .O(N__26980),
            .I(N__26977));
    LocalMux I__5603 (
            .O(N__26977),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__5602 (
            .O(N__26974),
            .I(N__26971));
    LocalMux I__5601 (
            .O(N__26971),
            .I(N__26968));
    Span4Mux_v I__5600 (
            .O(N__26968),
            .I(N__26965));
    Span4Mux_h I__5599 (
            .O(N__26965),
            .I(N__26962));
    Odrv4 I__5598 (
            .O(N__26962),
            .I(M_this_oam_ram_write_data_21));
    CascadeMux I__5597 (
            .O(N__26959),
            .I(N__26951));
    CascadeMux I__5596 (
            .O(N__26958),
            .I(N__26948));
    CascadeMux I__5595 (
            .O(N__26957),
            .I(N__26941));
    CascadeMux I__5594 (
            .O(N__26956),
            .I(N__26938));
    CascadeMux I__5593 (
            .O(N__26955),
            .I(N__26933));
    CascadeMux I__5592 (
            .O(N__26954),
            .I(N__26930));
    InMux I__5591 (
            .O(N__26951),
            .I(N__26927));
    InMux I__5590 (
            .O(N__26948),
            .I(N__26924));
    CascadeMux I__5589 (
            .O(N__26947),
            .I(N__26921));
    CascadeMux I__5588 (
            .O(N__26946),
            .I(N__26918));
    CascadeMux I__5587 (
            .O(N__26945),
            .I(N__26915));
    CascadeMux I__5586 (
            .O(N__26944),
            .I(N__26912));
    InMux I__5585 (
            .O(N__26941),
            .I(N__26908));
    InMux I__5584 (
            .O(N__26938),
            .I(N__26905));
    CascadeMux I__5583 (
            .O(N__26937),
            .I(N__26902));
    CascadeMux I__5582 (
            .O(N__26936),
            .I(N__26899));
    InMux I__5581 (
            .O(N__26933),
            .I(N__26894));
    InMux I__5580 (
            .O(N__26930),
            .I(N__26890));
    LocalMux I__5579 (
            .O(N__26927),
            .I(N__26885));
    LocalMux I__5578 (
            .O(N__26924),
            .I(N__26885));
    InMux I__5577 (
            .O(N__26921),
            .I(N__26882));
    InMux I__5576 (
            .O(N__26918),
            .I(N__26879));
    InMux I__5575 (
            .O(N__26915),
            .I(N__26876));
    InMux I__5574 (
            .O(N__26912),
            .I(N__26873));
    CascadeMux I__5573 (
            .O(N__26911),
            .I(N__26870));
    LocalMux I__5572 (
            .O(N__26908),
            .I(N__26865));
    LocalMux I__5571 (
            .O(N__26905),
            .I(N__26865));
    InMux I__5570 (
            .O(N__26902),
            .I(N__26862));
    InMux I__5569 (
            .O(N__26899),
            .I(N__26859));
    CascadeMux I__5568 (
            .O(N__26898),
            .I(N__26856));
    CascadeMux I__5567 (
            .O(N__26897),
            .I(N__26853));
    LocalMux I__5566 (
            .O(N__26894),
            .I(N__26850));
    CascadeMux I__5565 (
            .O(N__26893),
            .I(N__26847));
    LocalMux I__5564 (
            .O(N__26890),
            .I(N__26844));
    Span4Mux_v I__5563 (
            .O(N__26885),
            .I(N__26837));
    LocalMux I__5562 (
            .O(N__26882),
            .I(N__26837));
    LocalMux I__5561 (
            .O(N__26879),
            .I(N__26837));
    LocalMux I__5560 (
            .O(N__26876),
            .I(N__26832));
    LocalMux I__5559 (
            .O(N__26873),
            .I(N__26832));
    InMux I__5558 (
            .O(N__26870),
            .I(N__26829));
    Span4Mux_v I__5557 (
            .O(N__26865),
            .I(N__26822));
    LocalMux I__5556 (
            .O(N__26862),
            .I(N__26822));
    LocalMux I__5555 (
            .O(N__26859),
            .I(N__26822));
    InMux I__5554 (
            .O(N__26856),
            .I(N__26819));
    InMux I__5553 (
            .O(N__26853),
            .I(N__26816));
    Span4Mux_h I__5552 (
            .O(N__26850),
            .I(N__26813));
    InMux I__5551 (
            .O(N__26847),
            .I(N__26810));
    Span4Mux_v I__5550 (
            .O(N__26844),
            .I(N__26805));
    Span4Mux_v I__5549 (
            .O(N__26837),
            .I(N__26805));
    Span4Mux_v I__5548 (
            .O(N__26832),
            .I(N__26800));
    LocalMux I__5547 (
            .O(N__26829),
            .I(N__26800));
    Span4Mux_v I__5546 (
            .O(N__26822),
            .I(N__26793));
    LocalMux I__5545 (
            .O(N__26819),
            .I(N__26793));
    LocalMux I__5544 (
            .O(N__26816),
            .I(N__26793));
    Span4Mux_h I__5543 (
            .O(N__26813),
            .I(N__26790));
    LocalMux I__5542 (
            .O(N__26810),
            .I(N__26787));
    Span4Mux_h I__5541 (
            .O(N__26805),
            .I(N__26784));
    Span4Mux_v I__5540 (
            .O(N__26800),
            .I(N__26781));
    Span4Mux_v I__5539 (
            .O(N__26793),
            .I(N__26778));
    Span4Mux_h I__5538 (
            .O(N__26790),
            .I(N__26773));
    Span4Mux_h I__5537 (
            .O(N__26787),
            .I(N__26773));
    Span4Mux_h I__5536 (
            .O(N__26784),
            .I(N__26769));
    Span4Mux_h I__5535 (
            .O(N__26781),
            .I(N__26764));
    Span4Mux_h I__5534 (
            .O(N__26778),
            .I(N__26764));
    Span4Mux_h I__5533 (
            .O(N__26773),
            .I(N__26761));
    InMux I__5532 (
            .O(N__26772),
            .I(N__26758));
    Odrv4 I__5531 (
            .O(N__26769),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv4 I__5530 (
            .O(N__26764),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv4 I__5529 (
            .O(N__26761),
            .I(M_this_spr_address_qZ0Z_0));
    LocalMux I__5528 (
            .O(N__26758),
            .I(M_this_spr_address_qZ0Z_0));
    CascadeMux I__5527 (
            .O(N__26749),
            .I(N__26742));
    CascadeMux I__5526 (
            .O(N__26748),
            .I(N__26737));
    CascadeMux I__5525 (
            .O(N__26747),
            .I(N__26732));
    CascadeMux I__5524 (
            .O(N__26746),
            .I(N__26727));
    CascadeMux I__5523 (
            .O(N__26745),
            .I(N__26722));
    InMux I__5522 (
            .O(N__26742),
            .I(N__26718));
    CascadeMux I__5521 (
            .O(N__26741),
            .I(N__26715));
    CascadeMux I__5520 (
            .O(N__26740),
            .I(N__26712));
    InMux I__5519 (
            .O(N__26737),
            .I(N__26709));
    CascadeMux I__5518 (
            .O(N__26736),
            .I(N__26706));
    CascadeMux I__5517 (
            .O(N__26735),
            .I(N__26703));
    InMux I__5516 (
            .O(N__26732),
            .I(N__26700));
    CascadeMux I__5515 (
            .O(N__26731),
            .I(N__26697));
    CascadeMux I__5514 (
            .O(N__26730),
            .I(N__26694));
    InMux I__5513 (
            .O(N__26727),
            .I(N__26691));
    CascadeMux I__5512 (
            .O(N__26726),
            .I(N__26688));
    CascadeMux I__5511 (
            .O(N__26725),
            .I(N__26685));
    InMux I__5510 (
            .O(N__26722),
            .I(N__26682));
    CascadeMux I__5509 (
            .O(N__26721),
            .I(N__26679));
    LocalMux I__5508 (
            .O(N__26718),
            .I(N__26676));
    InMux I__5507 (
            .O(N__26715),
            .I(N__26673));
    InMux I__5506 (
            .O(N__26712),
            .I(N__26668));
    LocalMux I__5505 (
            .O(N__26709),
            .I(N__26665));
    InMux I__5504 (
            .O(N__26706),
            .I(N__26662));
    InMux I__5503 (
            .O(N__26703),
            .I(N__26659));
    LocalMux I__5502 (
            .O(N__26700),
            .I(N__26656));
    InMux I__5501 (
            .O(N__26697),
            .I(N__26653));
    InMux I__5500 (
            .O(N__26694),
            .I(N__26650));
    LocalMux I__5499 (
            .O(N__26691),
            .I(N__26647));
    InMux I__5498 (
            .O(N__26688),
            .I(N__26644));
    InMux I__5497 (
            .O(N__26685),
            .I(N__26641));
    LocalMux I__5496 (
            .O(N__26682),
            .I(N__26638));
    InMux I__5495 (
            .O(N__26679),
            .I(N__26635));
    Span4Mux_v I__5494 (
            .O(N__26676),
            .I(N__26630));
    LocalMux I__5493 (
            .O(N__26673),
            .I(N__26630));
    CascadeMux I__5492 (
            .O(N__26672),
            .I(N__26627));
    CascadeMux I__5491 (
            .O(N__26671),
            .I(N__26624));
    LocalMux I__5490 (
            .O(N__26668),
            .I(N__26617));
    Span4Mux_v I__5489 (
            .O(N__26665),
            .I(N__26617));
    LocalMux I__5488 (
            .O(N__26662),
            .I(N__26617));
    LocalMux I__5487 (
            .O(N__26659),
            .I(N__26614));
    Span4Mux_h I__5486 (
            .O(N__26656),
            .I(N__26611));
    LocalMux I__5485 (
            .O(N__26653),
            .I(N__26608));
    LocalMux I__5484 (
            .O(N__26650),
            .I(N__26603));
    Span4Mux_v I__5483 (
            .O(N__26647),
            .I(N__26603));
    LocalMux I__5482 (
            .O(N__26644),
            .I(N__26596));
    LocalMux I__5481 (
            .O(N__26641),
            .I(N__26596));
    Span4Mux_v I__5480 (
            .O(N__26638),
            .I(N__26596));
    LocalMux I__5479 (
            .O(N__26635),
            .I(N__26591));
    Span4Mux_h I__5478 (
            .O(N__26630),
            .I(N__26591));
    InMux I__5477 (
            .O(N__26627),
            .I(N__26588));
    InMux I__5476 (
            .O(N__26624),
            .I(N__26585));
    Span4Mux_v I__5475 (
            .O(N__26617),
            .I(N__26580));
    Span4Mux_v I__5474 (
            .O(N__26614),
            .I(N__26580));
    Span4Mux_v I__5473 (
            .O(N__26611),
            .I(N__26577));
    Sp12to4 I__5472 (
            .O(N__26608),
            .I(N__26573));
    Span4Mux_v I__5471 (
            .O(N__26603),
            .I(N__26568));
    Span4Mux_v I__5470 (
            .O(N__26596),
            .I(N__26568));
    Sp12to4 I__5469 (
            .O(N__26591),
            .I(N__26565));
    LocalMux I__5468 (
            .O(N__26588),
            .I(N__26562));
    LocalMux I__5467 (
            .O(N__26585),
            .I(N__26557));
    Sp12to4 I__5466 (
            .O(N__26580),
            .I(N__26557));
    Span4Mux_h I__5465 (
            .O(N__26577),
            .I(N__26554));
    InMux I__5464 (
            .O(N__26576),
            .I(N__26551));
    Span12Mux_v I__5463 (
            .O(N__26573),
            .I(N__26544));
    Sp12to4 I__5462 (
            .O(N__26568),
            .I(N__26544));
    Span12Mux_v I__5461 (
            .O(N__26565),
            .I(N__26544));
    Span12Mux_h I__5460 (
            .O(N__26562),
            .I(N__26539));
    Span12Mux_h I__5459 (
            .O(N__26557),
            .I(N__26539));
    Span4Mux_h I__5458 (
            .O(N__26554),
            .I(N__26536));
    LocalMux I__5457 (
            .O(N__26551),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv12 I__5456 (
            .O(N__26544),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv12 I__5455 (
            .O(N__26539),
            .I(M_this_spr_address_qZ0Z_1));
    Odrv4 I__5454 (
            .O(N__26536),
            .I(M_this_spr_address_qZ0Z_1));
    InMux I__5453 (
            .O(N__26527),
            .I(un1_M_this_spr_address_q_cry_0));
    CascadeMux I__5452 (
            .O(N__26524),
            .I(N__26518));
    CascadeMux I__5451 (
            .O(N__26523),
            .I(N__26515));
    CascadeMux I__5450 (
            .O(N__26522),
            .I(N__26509));
    CascadeMux I__5449 (
            .O(N__26521),
            .I(N__26505));
    InMux I__5448 (
            .O(N__26518),
            .I(N__26502));
    InMux I__5447 (
            .O(N__26515),
            .I(N__26499));
    CascadeMux I__5446 (
            .O(N__26514),
            .I(N__26496));
    CascadeMux I__5445 (
            .O(N__26513),
            .I(N__26493));
    CascadeMux I__5444 (
            .O(N__26512),
            .I(N__26490));
    InMux I__5443 (
            .O(N__26509),
            .I(N__26486));
    CascadeMux I__5442 (
            .O(N__26508),
            .I(N__26483));
    InMux I__5441 (
            .O(N__26505),
            .I(N__26479));
    LocalMux I__5440 (
            .O(N__26502),
            .I(N__26474));
    LocalMux I__5439 (
            .O(N__26499),
            .I(N__26474));
    InMux I__5438 (
            .O(N__26496),
            .I(N__26471));
    InMux I__5437 (
            .O(N__26493),
            .I(N__26468));
    InMux I__5436 (
            .O(N__26490),
            .I(N__26460));
    CascadeMux I__5435 (
            .O(N__26489),
            .I(N__26457));
    LocalMux I__5434 (
            .O(N__26486),
            .I(N__26453));
    InMux I__5433 (
            .O(N__26483),
            .I(N__26450));
    CascadeMux I__5432 (
            .O(N__26482),
            .I(N__26447));
    LocalMux I__5431 (
            .O(N__26479),
            .I(N__26444));
    Span4Mux_v I__5430 (
            .O(N__26474),
            .I(N__26437));
    LocalMux I__5429 (
            .O(N__26471),
            .I(N__26437));
    LocalMux I__5428 (
            .O(N__26468),
            .I(N__26437));
    CascadeMux I__5427 (
            .O(N__26467),
            .I(N__26434));
    CascadeMux I__5426 (
            .O(N__26466),
            .I(N__26431));
    CascadeMux I__5425 (
            .O(N__26465),
            .I(N__26428));
    CascadeMux I__5424 (
            .O(N__26464),
            .I(N__26425));
    CascadeMux I__5423 (
            .O(N__26463),
            .I(N__26422));
    LocalMux I__5422 (
            .O(N__26460),
            .I(N__26419));
    InMux I__5421 (
            .O(N__26457),
            .I(N__26416));
    CascadeMux I__5420 (
            .O(N__26456),
            .I(N__26413));
    Span4Mux_h I__5419 (
            .O(N__26453),
            .I(N__26410));
    LocalMux I__5418 (
            .O(N__26450),
            .I(N__26407));
    InMux I__5417 (
            .O(N__26447),
            .I(N__26404));
    Span4Mux_v I__5416 (
            .O(N__26444),
            .I(N__26399));
    Span4Mux_v I__5415 (
            .O(N__26437),
            .I(N__26399));
    InMux I__5414 (
            .O(N__26434),
            .I(N__26396));
    InMux I__5413 (
            .O(N__26431),
            .I(N__26393));
    InMux I__5412 (
            .O(N__26428),
            .I(N__26390));
    InMux I__5411 (
            .O(N__26425),
            .I(N__26387));
    InMux I__5410 (
            .O(N__26422),
            .I(N__26384));
    Span4Mux_v I__5409 (
            .O(N__26419),
            .I(N__26379));
    LocalMux I__5408 (
            .O(N__26416),
            .I(N__26379));
    InMux I__5407 (
            .O(N__26413),
            .I(N__26376));
    Span4Mux_h I__5406 (
            .O(N__26410),
            .I(N__26373));
    Span4Mux_h I__5405 (
            .O(N__26407),
            .I(N__26370));
    LocalMux I__5404 (
            .O(N__26404),
            .I(N__26367));
    Span4Mux_h I__5403 (
            .O(N__26399),
            .I(N__26364));
    LocalMux I__5402 (
            .O(N__26396),
            .I(N__26357));
    LocalMux I__5401 (
            .O(N__26393),
            .I(N__26357));
    LocalMux I__5400 (
            .O(N__26390),
            .I(N__26357));
    LocalMux I__5399 (
            .O(N__26387),
            .I(N__26348));
    LocalMux I__5398 (
            .O(N__26384),
            .I(N__26348));
    Sp12to4 I__5397 (
            .O(N__26379),
            .I(N__26348));
    LocalMux I__5396 (
            .O(N__26376),
            .I(N__26348));
    Span4Mux_h I__5395 (
            .O(N__26373),
            .I(N__26341));
    Span4Mux_v I__5394 (
            .O(N__26370),
            .I(N__26341));
    Span4Mux_h I__5393 (
            .O(N__26367),
            .I(N__26341));
    Sp12to4 I__5392 (
            .O(N__26364),
            .I(N__26333));
    Span12Mux_v I__5391 (
            .O(N__26357),
            .I(N__26333));
    Span12Mux_v I__5390 (
            .O(N__26348),
            .I(N__26333));
    Span4Mux_h I__5389 (
            .O(N__26341),
            .I(N__26330));
    InMux I__5388 (
            .O(N__26340),
            .I(N__26327));
    Odrv12 I__5387 (
            .O(N__26333),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv4 I__5386 (
            .O(N__26330),
            .I(M_this_spr_address_qZ0Z_2));
    LocalMux I__5385 (
            .O(N__26327),
            .I(M_this_spr_address_qZ0Z_2));
    InMux I__5384 (
            .O(N__26320),
            .I(un1_M_this_spr_address_q_cry_1));
    CascadeMux I__5383 (
            .O(N__26317),
            .I(N__26313));
    CascadeMux I__5382 (
            .O(N__26316),
            .I(N__26309));
    InMux I__5381 (
            .O(N__26313),
            .I(N__26304));
    CascadeMux I__5380 (
            .O(N__26312),
            .I(N__26301));
    InMux I__5379 (
            .O(N__26309),
            .I(N__26294));
    CascadeMux I__5378 (
            .O(N__26308),
            .I(N__26291));
    CascadeMux I__5377 (
            .O(N__26307),
            .I(N__26288));
    LocalMux I__5376 (
            .O(N__26304),
            .I(N__26285));
    InMux I__5375 (
            .O(N__26301),
            .I(N__26282));
    CascadeMux I__5374 (
            .O(N__26300),
            .I(N__26279));
    CascadeMux I__5373 (
            .O(N__26299),
            .I(N__26275));
    CascadeMux I__5372 (
            .O(N__26298),
            .I(N__26271));
    CascadeMux I__5371 (
            .O(N__26297),
            .I(N__26268));
    LocalMux I__5370 (
            .O(N__26294),
            .I(N__26265));
    InMux I__5369 (
            .O(N__26291),
            .I(N__26262));
    InMux I__5368 (
            .O(N__26288),
            .I(N__26258));
    Span4Mux_h I__5367 (
            .O(N__26285),
            .I(N__26255));
    LocalMux I__5366 (
            .O(N__26282),
            .I(N__26252));
    InMux I__5365 (
            .O(N__26279),
            .I(N__26249));
    CascadeMux I__5364 (
            .O(N__26278),
            .I(N__26246));
    InMux I__5363 (
            .O(N__26275),
            .I(N__26243));
    CascadeMux I__5362 (
            .O(N__26274),
            .I(N__26240));
    InMux I__5361 (
            .O(N__26271),
            .I(N__26236));
    InMux I__5360 (
            .O(N__26268),
            .I(N__26232));
    Span4Mux_h I__5359 (
            .O(N__26265),
            .I(N__26228));
    LocalMux I__5358 (
            .O(N__26262),
            .I(N__26225));
    CascadeMux I__5357 (
            .O(N__26261),
            .I(N__26222));
    LocalMux I__5356 (
            .O(N__26258),
            .I(N__26219));
    Span4Mux_v I__5355 (
            .O(N__26255),
            .I(N__26213));
    Span4Mux_h I__5354 (
            .O(N__26252),
            .I(N__26213));
    LocalMux I__5353 (
            .O(N__26249),
            .I(N__26210));
    InMux I__5352 (
            .O(N__26246),
            .I(N__26207));
    LocalMux I__5351 (
            .O(N__26243),
            .I(N__26204));
    InMux I__5350 (
            .O(N__26240),
            .I(N__26201));
    CascadeMux I__5349 (
            .O(N__26239),
            .I(N__26198));
    LocalMux I__5348 (
            .O(N__26236),
            .I(N__26195));
    CascadeMux I__5347 (
            .O(N__26235),
            .I(N__26192));
    LocalMux I__5346 (
            .O(N__26232),
            .I(N__26189));
    CascadeMux I__5345 (
            .O(N__26231),
            .I(N__26186));
    Span4Mux_v I__5344 (
            .O(N__26228),
            .I(N__26181));
    Span4Mux_h I__5343 (
            .O(N__26225),
            .I(N__26181));
    InMux I__5342 (
            .O(N__26222),
            .I(N__26178));
    Span4Mux_h I__5341 (
            .O(N__26219),
            .I(N__26175));
    CascadeMux I__5340 (
            .O(N__26218),
            .I(N__26172));
    Span4Mux_v I__5339 (
            .O(N__26213),
            .I(N__26167));
    Span4Mux_h I__5338 (
            .O(N__26210),
            .I(N__26167));
    LocalMux I__5337 (
            .O(N__26207),
            .I(N__26164));
    Span4Mux_h I__5336 (
            .O(N__26204),
            .I(N__26161));
    LocalMux I__5335 (
            .O(N__26201),
            .I(N__26158));
    InMux I__5334 (
            .O(N__26198),
            .I(N__26155));
    Span4Mux_s3_v I__5333 (
            .O(N__26195),
            .I(N__26152));
    InMux I__5332 (
            .O(N__26192),
            .I(N__26149));
    Span4Mux_v I__5331 (
            .O(N__26189),
            .I(N__26146));
    InMux I__5330 (
            .O(N__26186),
            .I(N__26143));
    Span4Mux_v I__5329 (
            .O(N__26181),
            .I(N__26138));
    LocalMux I__5328 (
            .O(N__26178),
            .I(N__26138));
    Span4Mux_v I__5327 (
            .O(N__26175),
            .I(N__26135));
    InMux I__5326 (
            .O(N__26172),
            .I(N__26132));
    Span4Mux_h I__5325 (
            .O(N__26167),
            .I(N__26129));
    Span4Mux_h I__5324 (
            .O(N__26164),
            .I(N__26126));
    Span4Mux_v I__5323 (
            .O(N__26161),
            .I(N__26121));
    Span4Mux_h I__5322 (
            .O(N__26158),
            .I(N__26121));
    LocalMux I__5321 (
            .O(N__26155),
            .I(N__26118));
    Sp12to4 I__5320 (
            .O(N__26152),
            .I(N__26113));
    LocalMux I__5319 (
            .O(N__26149),
            .I(N__26113));
    Sp12to4 I__5318 (
            .O(N__26146),
            .I(N__26108));
    LocalMux I__5317 (
            .O(N__26143),
            .I(N__26108));
    Sp12to4 I__5316 (
            .O(N__26138),
            .I(N__26105));
    Sp12to4 I__5315 (
            .O(N__26135),
            .I(N__26100));
    LocalMux I__5314 (
            .O(N__26132),
            .I(N__26100));
    Span4Mux_h I__5313 (
            .O(N__26129),
            .I(N__26091));
    Span4Mux_v I__5312 (
            .O(N__26126),
            .I(N__26091));
    Span4Mux_v I__5311 (
            .O(N__26121),
            .I(N__26091));
    Span4Mux_h I__5310 (
            .O(N__26118),
            .I(N__26091));
    Span12Mux_h I__5309 (
            .O(N__26113),
            .I(N__26085));
    Span12Mux_h I__5308 (
            .O(N__26108),
            .I(N__26085));
    Span12Mux_h I__5307 (
            .O(N__26105),
            .I(N__26080));
    Span12Mux_h I__5306 (
            .O(N__26100),
            .I(N__26080));
    Span4Mux_h I__5305 (
            .O(N__26091),
            .I(N__26077));
    InMux I__5304 (
            .O(N__26090),
            .I(N__26074));
    Odrv12 I__5303 (
            .O(N__26085),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv12 I__5302 (
            .O(N__26080),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv4 I__5301 (
            .O(N__26077),
            .I(M_this_spr_address_qZ0Z_3));
    LocalMux I__5300 (
            .O(N__26074),
            .I(M_this_spr_address_qZ0Z_3));
    InMux I__5299 (
            .O(N__26065),
            .I(un1_M_this_spr_address_q_cry_2));
    CascadeMux I__5298 (
            .O(N__26062),
            .I(N__26056));
    CascadeMux I__5297 (
            .O(N__26061),
            .I(N__26053));
    CascadeMux I__5296 (
            .O(N__26060),
            .I(N__26046));
    CascadeMux I__5295 (
            .O(N__26059),
            .I(N__26043));
    InMux I__5294 (
            .O(N__26056),
            .I(N__26036));
    InMux I__5293 (
            .O(N__26053),
            .I(N__26033));
    CascadeMux I__5292 (
            .O(N__26052),
            .I(N__26030));
    CascadeMux I__5291 (
            .O(N__26051),
            .I(N__26027));
    CascadeMux I__5290 (
            .O(N__26050),
            .I(N__26024));
    CascadeMux I__5289 (
            .O(N__26049),
            .I(N__26021));
    InMux I__5288 (
            .O(N__26046),
            .I(N__26018));
    InMux I__5287 (
            .O(N__26043),
            .I(N__26015));
    CascadeMux I__5286 (
            .O(N__26042),
            .I(N__26012));
    CascadeMux I__5285 (
            .O(N__26041),
            .I(N__26009));
    CascadeMux I__5284 (
            .O(N__26040),
            .I(N__26004));
    CascadeMux I__5283 (
            .O(N__26039),
            .I(N__26001));
    LocalMux I__5282 (
            .O(N__26036),
            .I(N__25994));
    LocalMux I__5281 (
            .O(N__26033),
            .I(N__25994));
    InMux I__5280 (
            .O(N__26030),
            .I(N__25991));
    InMux I__5279 (
            .O(N__26027),
            .I(N__25988));
    InMux I__5278 (
            .O(N__26024),
            .I(N__25985));
    InMux I__5277 (
            .O(N__26021),
            .I(N__25982));
    LocalMux I__5276 (
            .O(N__26018),
            .I(N__25977));
    LocalMux I__5275 (
            .O(N__26015),
            .I(N__25977));
    InMux I__5274 (
            .O(N__26012),
            .I(N__25974));
    InMux I__5273 (
            .O(N__26009),
            .I(N__25971));
    CascadeMux I__5272 (
            .O(N__26008),
            .I(N__25968));
    CascadeMux I__5271 (
            .O(N__26007),
            .I(N__25965));
    InMux I__5270 (
            .O(N__26004),
            .I(N__25962));
    InMux I__5269 (
            .O(N__26001),
            .I(N__25959));
    CascadeMux I__5268 (
            .O(N__26000),
            .I(N__25956));
    CascadeMux I__5267 (
            .O(N__25999),
            .I(N__25953));
    Span4Mux_v I__5266 (
            .O(N__25994),
            .I(N__25946));
    LocalMux I__5265 (
            .O(N__25991),
            .I(N__25946));
    LocalMux I__5264 (
            .O(N__25988),
            .I(N__25946));
    LocalMux I__5263 (
            .O(N__25985),
            .I(N__25941));
    LocalMux I__5262 (
            .O(N__25982),
            .I(N__25941));
    Span4Mux_v I__5261 (
            .O(N__25977),
            .I(N__25934));
    LocalMux I__5260 (
            .O(N__25974),
            .I(N__25934));
    LocalMux I__5259 (
            .O(N__25971),
            .I(N__25934));
    InMux I__5258 (
            .O(N__25968),
            .I(N__25931));
    InMux I__5257 (
            .O(N__25965),
            .I(N__25928));
    LocalMux I__5256 (
            .O(N__25962),
            .I(N__25923));
    LocalMux I__5255 (
            .O(N__25959),
            .I(N__25923));
    InMux I__5254 (
            .O(N__25956),
            .I(N__25920));
    InMux I__5253 (
            .O(N__25953),
            .I(N__25917));
    Span4Mux_v I__5252 (
            .O(N__25946),
            .I(N__25912));
    Span4Mux_v I__5251 (
            .O(N__25941),
            .I(N__25912));
    Span4Mux_v I__5250 (
            .O(N__25934),
            .I(N__25905));
    LocalMux I__5249 (
            .O(N__25931),
            .I(N__25905));
    LocalMux I__5248 (
            .O(N__25928),
            .I(N__25905));
    Span4Mux_v I__5247 (
            .O(N__25923),
            .I(N__25898));
    LocalMux I__5246 (
            .O(N__25920),
            .I(N__25898));
    LocalMux I__5245 (
            .O(N__25917),
            .I(N__25898));
    Span4Mux_h I__5244 (
            .O(N__25912),
            .I(N__25895));
    Span4Mux_v I__5243 (
            .O(N__25905),
            .I(N__25890));
    Span4Mux_v I__5242 (
            .O(N__25898),
            .I(N__25890));
    Span4Mux_h I__5241 (
            .O(N__25895),
            .I(N__25884));
    Span4Mux_h I__5240 (
            .O(N__25890),
            .I(N__25884));
    InMux I__5239 (
            .O(N__25889),
            .I(N__25881));
    Odrv4 I__5238 (
            .O(N__25884),
            .I(M_this_spr_address_qZ0Z_4));
    LocalMux I__5237 (
            .O(N__25881),
            .I(M_this_spr_address_qZ0Z_4));
    InMux I__5236 (
            .O(N__25876),
            .I(un1_M_this_spr_address_q_cry_3));
    CascadeMux I__5235 (
            .O(N__25873),
            .I(N__25870));
    InMux I__5234 (
            .O(N__25870),
            .I(N__25861));
    CascadeMux I__5233 (
            .O(N__25869),
            .I(N__25858));
    CascadeMux I__5232 (
            .O(N__25868),
            .I(N__25854));
    CascadeMux I__5231 (
            .O(N__25867),
            .I(N__25850));
    CascadeMux I__5230 (
            .O(N__25866),
            .I(N__25847));
    CascadeMux I__5229 (
            .O(N__25865),
            .I(N__25844));
    CascadeMux I__5228 (
            .O(N__25864),
            .I(N__25837));
    LocalMux I__5227 (
            .O(N__25861),
            .I(N__25833));
    InMux I__5226 (
            .O(N__25858),
            .I(N__25830));
    CascadeMux I__5225 (
            .O(N__25857),
            .I(N__25827));
    InMux I__5224 (
            .O(N__25854),
            .I(N__25824));
    CascadeMux I__5223 (
            .O(N__25853),
            .I(N__25821));
    InMux I__5222 (
            .O(N__25850),
            .I(N__25818));
    InMux I__5221 (
            .O(N__25847),
            .I(N__25815));
    InMux I__5220 (
            .O(N__25844),
            .I(N__25812));
    CascadeMux I__5219 (
            .O(N__25843),
            .I(N__25809));
    CascadeMux I__5218 (
            .O(N__25842),
            .I(N__25806));
    CascadeMux I__5217 (
            .O(N__25841),
            .I(N__25803));
    CascadeMux I__5216 (
            .O(N__25840),
            .I(N__25800));
    InMux I__5215 (
            .O(N__25837),
            .I(N__25797));
    CascadeMux I__5214 (
            .O(N__25836),
            .I(N__25794));
    Span4Mux_v I__5213 (
            .O(N__25833),
            .I(N__25787));
    LocalMux I__5212 (
            .O(N__25830),
            .I(N__25787));
    InMux I__5211 (
            .O(N__25827),
            .I(N__25784));
    LocalMux I__5210 (
            .O(N__25824),
            .I(N__25781));
    InMux I__5209 (
            .O(N__25821),
            .I(N__25778));
    LocalMux I__5208 (
            .O(N__25818),
            .I(N__25775));
    LocalMux I__5207 (
            .O(N__25815),
            .I(N__25770));
    LocalMux I__5206 (
            .O(N__25812),
            .I(N__25770));
    InMux I__5205 (
            .O(N__25809),
            .I(N__25767));
    InMux I__5204 (
            .O(N__25806),
            .I(N__25764));
    InMux I__5203 (
            .O(N__25803),
            .I(N__25761));
    InMux I__5202 (
            .O(N__25800),
            .I(N__25758));
    LocalMux I__5201 (
            .O(N__25797),
            .I(N__25755));
    InMux I__5200 (
            .O(N__25794),
            .I(N__25752));
    CascadeMux I__5199 (
            .O(N__25793),
            .I(N__25749));
    CascadeMux I__5198 (
            .O(N__25792),
            .I(N__25746));
    Span4Mux_v I__5197 (
            .O(N__25787),
            .I(N__25743));
    LocalMux I__5196 (
            .O(N__25784),
            .I(N__25736));
    Span4Mux_v I__5195 (
            .O(N__25781),
            .I(N__25736));
    LocalMux I__5194 (
            .O(N__25778),
            .I(N__25736));
    Span4Mux_s3_v I__5193 (
            .O(N__25775),
            .I(N__25733));
    Span4Mux_v I__5192 (
            .O(N__25770),
            .I(N__25728));
    LocalMux I__5191 (
            .O(N__25767),
            .I(N__25728));
    LocalMux I__5190 (
            .O(N__25764),
            .I(N__25723));
    LocalMux I__5189 (
            .O(N__25761),
            .I(N__25723));
    LocalMux I__5188 (
            .O(N__25758),
            .I(N__25720));
    Span4Mux_h I__5187 (
            .O(N__25755),
            .I(N__25717));
    LocalMux I__5186 (
            .O(N__25752),
            .I(N__25714));
    InMux I__5185 (
            .O(N__25749),
            .I(N__25711));
    InMux I__5184 (
            .O(N__25746),
            .I(N__25708));
    Span4Mux_v I__5183 (
            .O(N__25743),
            .I(N__25703));
    Span4Mux_v I__5182 (
            .O(N__25736),
            .I(N__25703));
    Span4Mux_h I__5181 (
            .O(N__25733),
            .I(N__25698));
    Span4Mux_h I__5180 (
            .O(N__25728),
            .I(N__25698));
    Span4Mux_v I__5179 (
            .O(N__25723),
            .I(N__25693));
    Span4Mux_v I__5178 (
            .O(N__25720),
            .I(N__25693));
    Span4Mux_v I__5177 (
            .O(N__25717),
            .I(N__25688));
    Span4Mux_h I__5176 (
            .O(N__25714),
            .I(N__25688));
    LocalMux I__5175 (
            .O(N__25711),
            .I(N__25684));
    LocalMux I__5174 (
            .O(N__25708),
            .I(N__25679));
    Sp12to4 I__5173 (
            .O(N__25703),
            .I(N__25679));
    Sp12to4 I__5172 (
            .O(N__25698),
            .I(N__25676));
    Span4Mux_h I__5171 (
            .O(N__25693),
            .I(N__25673));
    Span4Mux_h I__5170 (
            .O(N__25688),
            .I(N__25670));
    InMux I__5169 (
            .O(N__25687),
            .I(N__25667));
    Span12Mux_h I__5168 (
            .O(N__25684),
            .I(N__25662));
    Span12Mux_h I__5167 (
            .O(N__25679),
            .I(N__25662));
    Span12Mux_v I__5166 (
            .O(N__25676),
            .I(N__25659));
    Odrv4 I__5165 (
            .O(N__25673),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv4 I__5164 (
            .O(N__25670),
            .I(M_this_spr_address_qZ0Z_5));
    LocalMux I__5163 (
            .O(N__25667),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv12 I__5162 (
            .O(N__25662),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv12 I__5161 (
            .O(N__25659),
            .I(M_this_spr_address_qZ0Z_5));
    InMux I__5160 (
            .O(N__25648),
            .I(un1_M_this_spr_address_q_cry_4));
    CascadeMux I__5159 (
            .O(N__25645),
            .I(N__25642));
    InMux I__5158 (
            .O(N__25642),
            .I(N__25634));
    CascadeMux I__5157 (
            .O(N__25641),
            .I(N__25631));
    CascadeMux I__5156 (
            .O(N__25640),
            .I(N__25627));
    CascadeMux I__5155 (
            .O(N__25639),
            .I(N__25623));
    CascadeMux I__5154 (
            .O(N__25638),
            .I(N__25620));
    CascadeMux I__5153 (
            .O(N__25637),
            .I(N__25615));
    LocalMux I__5152 (
            .O(N__25634),
            .I(N__25611));
    InMux I__5151 (
            .O(N__25631),
            .I(N__25608));
    CascadeMux I__5150 (
            .O(N__25630),
            .I(N__25605));
    InMux I__5149 (
            .O(N__25627),
            .I(N__25601));
    CascadeMux I__5148 (
            .O(N__25626),
            .I(N__25598));
    InMux I__5147 (
            .O(N__25623),
            .I(N__25594));
    InMux I__5146 (
            .O(N__25620),
            .I(N__25591));
    CascadeMux I__5145 (
            .O(N__25619),
            .I(N__25588));
    CascadeMux I__5144 (
            .O(N__25618),
            .I(N__25585));
    InMux I__5143 (
            .O(N__25615),
            .I(N__25581));
    CascadeMux I__5142 (
            .O(N__25614),
            .I(N__25578));
    Span4Mux_h I__5141 (
            .O(N__25611),
            .I(N__25574));
    LocalMux I__5140 (
            .O(N__25608),
            .I(N__25571));
    InMux I__5139 (
            .O(N__25605),
            .I(N__25568));
    CascadeMux I__5138 (
            .O(N__25604),
            .I(N__25565));
    LocalMux I__5137 (
            .O(N__25601),
            .I(N__25562));
    InMux I__5136 (
            .O(N__25598),
            .I(N__25559));
    CascadeMux I__5135 (
            .O(N__25597),
            .I(N__25556));
    LocalMux I__5134 (
            .O(N__25594),
            .I(N__25552));
    LocalMux I__5133 (
            .O(N__25591),
            .I(N__25549));
    InMux I__5132 (
            .O(N__25588),
            .I(N__25546));
    InMux I__5131 (
            .O(N__25585),
            .I(N__25543));
    CascadeMux I__5130 (
            .O(N__25584),
            .I(N__25540));
    LocalMux I__5129 (
            .O(N__25581),
            .I(N__25537));
    InMux I__5128 (
            .O(N__25578),
            .I(N__25534));
    CascadeMux I__5127 (
            .O(N__25577),
            .I(N__25531));
    Span4Mux_v I__5126 (
            .O(N__25574),
            .I(N__25526));
    Span4Mux_h I__5125 (
            .O(N__25571),
            .I(N__25526));
    LocalMux I__5124 (
            .O(N__25568),
            .I(N__25523));
    InMux I__5123 (
            .O(N__25565),
            .I(N__25520));
    Span4Mux_h I__5122 (
            .O(N__25562),
            .I(N__25517));
    LocalMux I__5121 (
            .O(N__25559),
            .I(N__25514));
    InMux I__5120 (
            .O(N__25556),
            .I(N__25511));
    CascadeMux I__5119 (
            .O(N__25555),
            .I(N__25508));
    Span4Mux_h I__5118 (
            .O(N__25552),
            .I(N__25505));
    Span4Mux_h I__5117 (
            .O(N__25549),
            .I(N__25502));
    LocalMux I__5116 (
            .O(N__25546),
            .I(N__25499));
    LocalMux I__5115 (
            .O(N__25543),
            .I(N__25496));
    InMux I__5114 (
            .O(N__25540),
            .I(N__25493));
    Span4Mux_h I__5113 (
            .O(N__25537),
            .I(N__25490));
    LocalMux I__5112 (
            .O(N__25534),
            .I(N__25487));
    InMux I__5111 (
            .O(N__25531),
            .I(N__25484));
    Span4Mux_v I__5110 (
            .O(N__25526),
            .I(N__25479));
    Span4Mux_h I__5109 (
            .O(N__25523),
            .I(N__25479));
    LocalMux I__5108 (
            .O(N__25520),
            .I(N__25476));
    Span4Mux_v I__5107 (
            .O(N__25517),
            .I(N__25471));
    Span4Mux_h I__5106 (
            .O(N__25514),
            .I(N__25471));
    LocalMux I__5105 (
            .O(N__25511),
            .I(N__25468));
    InMux I__5104 (
            .O(N__25508),
            .I(N__25465));
    Span4Mux_v I__5103 (
            .O(N__25505),
            .I(N__25458));
    Span4Mux_v I__5102 (
            .O(N__25502),
            .I(N__25458));
    Span4Mux_h I__5101 (
            .O(N__25499),
            .I(N__25458));
    Span4Mux_h I__5100 (
            .O(N__25496),
            .I(N__25455));
    LocalMux I__5099 (
            .O(N__25493),
            .I(N__25452));
    Span4Mux_v I__5098 (
            .O(N__25490),
            .I(N__25447));
    Span4Mux_h I__5097 (
            .O(N__25487),
            .I(N__25447));
    LocalMux I__5096 (
            .O(N__25484),
            .I(N__25444));
    Span4Mux_h I__5095 (
            .O(N__25479),
            .I(N__25441));
    Span4Mux_h I__5094 (
            .O(N__25476),
            .I(N__25438));
    Span4Mux_v I__5093 (
            .O(N__25471),
            .I(N__25433));
    Span4Mux_h I__5092 (
            .O(N__25468),
            .I(N__25433));
    LocalMux I__5091 (
            .O(N__25465),
            .I(N__25430));
    Span4Mux_h I__5090 (
            .O(N__25458),
            .I(N__25427));
    Span4Mux_v I__5089 (
            .O(N__25455),
            .I(N__25422));
    Span4Mux_h I__5088 (
            .O(N__25452),
            .I(N__25422));
    Span4Mux_v I__5087 (
            .O(N__25447),
            .I(N__25417));
    Span4Mux_h I__5086 (
            .O(N__25444),
            .I(N__25417));
    Span4Mux_h I__5085 (
            .O(N__25441),
            .I(N__25408));
    Span4Mux_v I__5084 (
            .O(N__25438),
            .I(N__25408));
    Span4Mux_v I__5083 (
            .O(N__25433),
            .I(N__25408));
    Span4Mux_h I__5082 (
            .O(N__25430),
            .I(N__25408));
    Span4Mux_h I__5081 (
            .O(N__25427),
            .I(N__25400));
    Span4Mux_h I__5080 (
            .O(N__25422),
            .I(N__25400));
    Span4Mux_h I__5079 (
            .O(N__25417),
            .I(N__25400));
    Span4Mux_h I__5078 (
            .O(N__25408),
            .I(N__25397));
    InMux I__5077 (
            .O(N__25407),
            .I(N__25394));
    Odrv4 I__5076 (
            .O(N__25400),
            .I(M_this_spr_address_qZ0Z_6));
    Odrv4 I__5075 (
            .O(N__25397),
            .I(M_this_spr_address_qZ0Z_6));
    LocalMux I__5074 (
            .O(N__25394),
            .I(M_this_spr_address_qZ0Z_6));
    InMux I__5073 (
            .O(N__25387),
            .I(un1_M_this_spr_address_q_cry_5));
    CascadeMux I__5072 (
            .O(N__25384),
            .I(N__25381));
    CascadeBuf I__5071 (
            .O(N__25381),
            .I(N__25378));
    CascadeMux I__5070 (
            .O(N__25378),
            .I(N__25374));
    CascadeMux I__5069 (
            .O(N__25377),
            .I(N__25371));
    InMux I__5068 (
            .O(N__25374),
            .I(N__25368));
    InMux I__5067 (
            .O(N__25371),
            .I(N__25363));
    LocalMux I__5066 (
            .O(N__25368),
            .I(N__25360));
    InMux I__5065 (
            .O(N__25367),
            .I(N__25357));
    InMux I__5064 (
            .O(N__25366),
            .I(N__25354));
    LocalMux I__5063 (
            .O(N__25363),
            .I(N__25351));
    Span12Mux_h I__5062 (
            .O(N__25360),
            .I(N__25348));
    LocalMux I__5061 (
            .O(N__25357),
            .I(M_this_ppu_oam_addr_4));
    LocalMux I__5060 (
            .O(N__25354),
            .I(M_this_ppu_oam_addr_4));
    Odrv4 I__5059 (
            .O(N__25351),
            .I(M_this_ppu_oam_addr_4));
    Odrv12 I__5058 (
            .O(N__25348),
            .I(M_this_ppu_oam_addr_4));
    InMux I__5057 (
            .O(N__25339),
            .I(N__25336));
    LocalMux I__5056 (
            .O(N__25336),
            .I(N__25333));
    Span4Mux_v I__5055 (
            .O(N__25333),
            .I(N__25330));
    Odrv4 I__5054 (
            .O(N__25330),
            .I(M_this_data_tmp_qZ0Z_13));
    InMux I__5053 (
            .O(N__25327),
            .I(N__25324));
    LocalMux I__5052 (
            .O(N__25324),
            .I(N__25321));
    Span4Mux_v I__5051 (
            .O(N__25321),
            .I(N__25318));
    Span4Mux_h I__5050 (
            .O(N__25318),
            .I(N__25315));
    Odrv4 I__5049 (
            .O(N__25315),
            .I(M_this_oam_ram_write_data_13));
    CascadeMux I__5048 (
            .O(N__25312),
            .I(N__25309));
    CascadeBuf I__5047 (
            .O(N__25309),
            .I(N__25306));
    CascadeMux I__5046 (
            .O(N__25306),
            .I(N__25303));
    InMux I__5045 (
            .O(N__25303),
            .I(N__25300));
    LocalMux I__5044 (
            .O(N__25300),
            .I(N__25297));
    Span4Mux_v I__5043 (
            .O(N__25297),
            .I(N__25291));
    InMux I__5042 (
            .O(N__25296),
            .I(N__25288));
    InMux I__5041 (
            .O(N__25295),
            .I(N__25285));
    InMux I__5040 (
            .O(N__25294),
            .I(N__25282));
    Span4Mux_h I__5039 (
            .O(N__25291),
            .I(N__25279));
    LocalMux I__5038 (
            .O(N__25288),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__5037 (
            .O(N__25285),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__5036 (
            .O(N__25282),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv4 I__5035 (
            .O(N__25279),
            .I(M_this_oam_address_qZ0Z_2));
    CascadeMux I__5034 (
            .O(N__25270),
            .I(N__25267));
    CascadeBuf I__5033 (
            .O(N__25267),
            .I(N__25264));
    CascadeMux I__5032 (
            .O(N__25264),
            .I(N__25261));
    InMux I__5031 (
            .O(N__25261),
            .I(N__25258));
    LocalMux I__5030 (
            .O(N__25258),
            .I(N__25255));
    Span4Mux_v I__5029 (
            .O(N__25255),
            .I(N__25251));
    CascadeMux I__5028 (
            .O(N__25254),
            .I(N__25248));
    Span4Mux_h I__5027 (
            .O(N__25251),
            .I(N__25244));
    InMux I__5026 (
            .O(N__25248),
            .I(N__25241));
    InMux I__5025 (
            .O(N__25247),
            .I(N__25238));
    Span4Mux_v I__5024 (
            .O(N__25244),
            .I(N__25235));
    LocalMux I__5023 (
            .O(N__25241),
            .I(M_this_oam_address_qZ0Z_3));
    LocalMux I__5022 (
            .O(N__25238),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv4 I__5021 (
            .O(N__25235),
            .I(M_this_oam_address_qZ0Z_3));
    InMux I__5020 (
            .O(N__25228),
            .I(N__25224));
    InMux I__5019 (
            .O(N__25227),
            .I(N__25221));
    LocalMux I__5018 (
            .O(N__25224),
            .I(N__25215));
    LocalMux I__5017 (
            .O(N__25221),
            .I(N__25215));
    InMux I__5016 (
            .O(N__25220),
            .I(N__25212));
    Sp12to4 I__5015 (
            .O(N__25215),
            .I(N__25207));
    LocalMux I__5014 (
            .O(N__25212),
            .I(N__25207));
    Odrv12 I__5013 (
            .O(N__25207),
            .I(un1_M_this_oam_address_q_c2));
    InMux I__5012 (
            .O(N__25204),
            .I(N__25198));
    InMux I__5011 (
            .O(N__25203),
            .I(N__25198));
    LocalMux I__5010 (
            .O(N__25198),
            .I(un1_M_this_oam_address_q_c4));
    CascadeMux I__5009 (
            .O(N__25195),
            .I(N__25192));
    CascadeBuf I__5008 (
            .O(N__25192),
            .I(N__25189));
    CascadeMux I__5007 (
            .O(N__25189),
            .I(N__25186));
    InMux I__5006 (
            .O(N__25186),
            .I(N__25183));
    LocalMux I__5005 (
            .O(N__25183),
            .I(N__25180));
    Span4Mux_v I__5004 (
            .O(N__25180),
            .I(N__25175));
    CascadeMux I__5003 (
            .O(N__25179),
            .I(N__25172));
    InMux I__5002 (
            .O(N__25178),
            .I(N__25169));
    Span4Mux_h I__5001 (
            .O(N__25175),
            .I(N__25166));
    InMux I__5000 (
            .O(N__25172),
            .I(N__25163));
    LocalMux I__4999 (
            .O(N__25169),
            .I(N__25158));
    Span4Mux_h I__4998 (
            .O(N__25166),
            .I(N__25158));
    LocalMux I__4997 (
            .O(N__25163),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__4996 (
            .O(N__25158),
            .I(M_this_oam_address_qZ0Z_5));
    CascadeMux I__4995 (
            .O(N__25153),
            .I(un1_M_this_oam_address_q_c4_cascade_));
    CascadeMux I__4994 (
            .O(N__25150),
            .I(N__25147));
    CascadeBuf I__4993 (
            .O(N__25147),
            .I(N__25144));
    CascadeMux I__4992 (
            .O(N__25144),
            .I(N__25141));
    InMux I__4991 (
            .O(N__25141),
            .I(N__25138));
    LocalMux I__4990 (
            .O(N__25138),
            .I(N__25135));
    Span4Mux_v I__4989 (
            .O(N__25135),
            .I(N__25132));
    Span4Mux_h I__4988 (
            .O(N__25132),
            .I(N__25126));
    InMux I__4987 (
            .O(N__25131),
            .I(N__25121));
    InMux I__4986 (
            .O(N__25130),
            .I(N__25121));
    InMux I__4985 (
            .O(N__25129),
            .I(N__25118));
    Span4Mux_h I__4984 (
            .O(N__25126),
            .I(N__25115));
    LocalMux I__4983 (
            .O(N__25121),
            .I(M_this_oam_address_qZ0Z_4));
    LocalMux I__4982 (
            .O(N__25118),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__4981 (
            .O(N__25115),
            .I(M_this_oam_address_qZ0Z_4));
    InMux I__4980 (
            .O(N__25108),
            .I(N__25104));
    InMux I__4979 (
            .O(N__25107),
            .I(N__25101));
    LocalMux I__4978 (
            .O(N__25104),
            .I(un1_M_this_oam_address_q_c6));
    LocalMux I__4977 (
            .O(N__25101),
            .I(un1_M_this_oam_address_q_c6));
    InMux I__4976 (
            .O(N__25096),
            .I(N__25086));
    InMux I__4975 (
            .O(N__25095),
            .I(N__25086));
    InMux I__4974 (
            .O(N__25094),
            .I(N__25081));
    InMux I__4973 (
            .O(N__25093),
            .I(N__25081));
    InMux I__4972 (
            .O(N__25092),
            .I(N__25078));
    InMux I__4971 (
            .O(N__25091),
            .I(N__25075));
    LocalMux I__4970 (
            .O(N__25086),
            .I(\this_ppu.N_268_i_0_0 ));
    LocalMux I__4969 (
            .O(N__25081),
            .I(\this_ppu.N_268_i_0_0 ));
    LocalMux I__4968 (
            .O(N__25078),
            .I(\this_ppu.N_268_i_0_0 ));
    LocalMux I__4967 (
            .O(N__25075),
            .I(\this_ppu.N_268_i_0_0 ));
    InMux I__4966 (
            .O(N__25066),
            .I(N__25052));
    InMux I__4965 (
            .O(N__25065),
            .I(N__25052));
    InMux I__4964 (
            .O(N__25064),
            .I(N__25052));
    InMux I__4963 (
            .O(N__25063),
            .I(N__25052));
    InMux I__4962 (
            .O(N__25062),
            .I(N__25049));
    InMux I__4961 (
            .O(N__25061),
            .I(N__25046));
    LocalMux I__4960 (
            .O(N__25052),
            .I(\this_ppu.N_1323_0 ));
    LocalMux I__4959 (
            .O(N__25049),
            .I(\this_ppu.N_1323_0 ));
    LocalMux I__4958 (
            .O(N__25046),
            .I(\this_ppu.N_1323_0 ));
    InMux I__4957 (
            .O(N__25039),
            .I(N__25035));
    InMux I__4956 (
            .O(N__25038),
            .I(N__25031));
    LocalMux I__4955 (
            .O(N__25035),
            .I(N__25028));
    InMux I__4954 (
            .O(N__25034),
            .I(N__25025));
    LocalMux I__4953 (
            .O(N__25031),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    Odrv4 I__4952 (
            .O(N__25028),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    LocalMux I__4951 (
            .O(N__25025),
            .I(\this_ppu.M_count_qZ0Z_0 ));
    CascadeMux I__4950 (
            .O(N__25018),
            .I(N__25015));
    InMux I__4949 (
            .O(N__25015),
            .I(N__25007));
    CascadeMux I__4948 (
            .O(N__25014),
            .I(N__25003));
    InMux I__4947 (
            .O(N__25013),
            .I(N__24998));
    InMux I__4946 (
            .O(N__25012),
            .I(N__24998));
    InMux I__4945 (
            .O(N__25011),
            .I(N__24995));
    CascadeMux I__4944 (
            .O(N__25010),
            .I(N__24990));
    LocalMux I__4943 (
            .O(N__25007),
            .I(N__24987));
    InMux I__4942 (
            .O(N__25006),
            .I(N__24984));
    InMux I__4941 (
            .O(N__25003),
            .I(N__24981));
    LocalMux I__4940 (
            .O(N__24998),
            .I(N__24976));
    LocalMux I__4939 (
            .O(N__24995),
            .I(N__24976));
    InMux I__4938 (
            .O(N__24994),
            .I(N__24969));
    InMux I__4937 (
            .O(N__24993),
            .I(N__24969));
    InMux I__4936 (
            .O(N__24990),
            .I(N__24969));
    Span4Mux_h I__4935 (
            .O(N__24987),
            .I(N__24966));
    LocalMux I__4934 (
            .O(N__24984),
            .I(N__24963));
    LocalMux I__4933 (
            .O(N__24981),
            .I(N__24956));
    Sp12to4 I__4932 (
            .O(N__24976),
            .I(N__24956));
    LocalMux I__4931 (
            .O(N__24969),
            .I(N__24956));
    Odrv4 I__4930 (
            .O(N__24966),
            .I(N_611));
    Odrv12 I__4929 (
            .O(N__24963),
            .I(N_611));
    Odrv12 I__4928 (
            .O(N__24956),
            .I(N_611));
    CascadeMux I__4927 (
            .O(N__24949),
            .I(N__24946));
    InMux I__4926 (
            .O(N__24946),
            .I(N__24943));
    LocalMux I__4925 (
            .O(N__24943),
            .I(N__24940));
    Odrv4 I__4924 (
            .O(N__24940),
            .I(M_this_data_count_q_s_13));
    CascadeMux I__4923 (
            .O(N__24937),
            .I(N__24934));
    InMux I__4922 (
            .O(N__24934),
            .I(N__24930));
    InMux I__4921 (
            .O(N__24933),
            .I(N__24927));
    LocalMux I__4920 (
            .O(N__24930),
            .I(N__24924));
    LocalMux I__4919 (
            .O(N__24927),
            .I(N__24919));
    Span4Mux_h I__4918 (
            .O(N__24924),
            .I(N__24919));
    Odrv4 I__4917 (
            .O(N__24919),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__4916 (
            .O(N__24916),
            .I(N__24913));
    LocalMux I__4915 (
            .O(N__24913),
            .I(M_this_data_count_q_s_8));
    CascadeMux I__4914 (
            .O(N__24910),
            .I(N__24905));
    InMux I__4913 (
            .O(N__24909),
            .I(N__24889));
    InMux I__4912 (
            .O(N__24908),
            .I(N__24889));
    InMux I__4911 (
            .O(N__24905),
            .I(N__24889));
    InMux I__4910 (
            .O(N__24904),
            .I(N__24889));
    InMux I__4909 (
            .O(N__24903),
            .I(N__24886));
    InMux I__4908 (
            .O(N__24902),
            .I(N__24877));
    InMux I__4907 (
            .O(N__24901),
            .I(N__24877));
    InMux I__4906 (
            .O(N__24900),
            .I(N__24877));
    InMux I__4905 (
            .O(N__24899),
            .I(N__24877));
    InMux I__4904 (
            .O(N__24898),
            .I(N__24870));
    LocalMux I__4903 (
            .O(N__24889),
            .I(N__24865));
    LocalMux I__4902 (
            .O(N__24886),
            .I(N__24865));
    LocalMux I__4901 (
            .O(N__24877),
            .I(N__24862));
    InMux I__4900 (
            .O(N__24876),
            .I(N__24853));
    InMux I__4899 (
            .O(N__24875),
            .I(N__24853));
    InMux I__4898 (
            .O(N__24874),
            .I(N__24853));
    InMux I__4897 (
            .O(N__24873),
            .I(N__24853));
    LocalMux I__4896 (
            .O(N__24870),
            .I(N__24850));
    Span4Mux_v I__4895 (
            .O(N__24865),
            .I(N__24847));
    Span4Mux_h I__4894 (
            .O(N__24862),
            .I(N__24842));
    LocalMux I__4893 (
            .O(N__24853),
            .I(N__24842));
    Odrv12 I__4892 (
            .O(N__24850),
            .I(N_660_i));
    Odrv4 I__4891 (
            .O(N__24847),
            .I(N_660_i));
    Odrv4 I__4890 (
            .O(N__24842),
            .I(N_660_i));
    InMux I__4889 (
            .O(N__24835),
            .I(N__24831));
    InMux I__4888 (
            .O(N__24834),
            .I(N__24828));
    LocalMux I__4887 (
            .O(N__24831),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__4886 (
            .O(N__24828),
            .I(M_this_data_count_qZ0Z_8));
    CEMux I__4885 (
            .O(N__24823),
            .I(N__24820));
    LocalMux I__4884 (
            .O(N__24820),
            .I(N__24816));
    CEMux I__4883 (
            .O(N__24819),
            .I(N__24812));
    Span4Mux_v I__4882 (
            .O(N__24816),
            .I(N__24808));
    CEMux I__4881 (
            .O(N__24815),
            .I(N__24805));
    LocalMux I__4880 (
            .O(N__24812),
            .I(N__24801));
    CEMux I__4879 (
            .O(N__24811),
            .I(N__24798));
    Span4Mux_h I__4878 (
            .O(N__24808),
            .I(N__24793));
    LocalMux I__4877 (
            .O(N__24805),
            .I(N__24793));
    CEMux I__4876 (
            .O(N__24804),
            .I(N__24790));
    Span4Mux_h I__4875 (
            .O(N__24801),
            .I(N__24785));
    LocalMux I__4874 (
            .O(N__24798),
            .I(N__24785));
    Span4Mux_v I__4873 (
            .O(N__24793),
            .I(N__24782));
    LocalMux I__4872 (
            .O(N__24790),
            .I(N__24779));
    Span4Mux_h I__4871 (
            .O(N__24785),
            .I(N__24776));
    Odrv4 I__4870 (
            .O(N__24782),
            .I(N_257));
    Odrv12 I__4869 (
            .O(N__24779),
            .I(N_257));
    Odrv4 I__4868 (
            .O(N__24776),
            .I(N_257));
    InMux I__4867 (
            .O(N__24769),
            .I(N__24766));
    LocalMux I__4866 (
            .O(N__24766),
            .I(N__24761));
    InMux I__4865 (
            .O(N__24765),
            .I(N__24758));
    InMux I__4864 (
            .O(N__24764),
            .I(N__24754));
    Span4Mux_v I__4863 (
            .O(N__24761),
            .I(N__24749));
    LocalMux I__4862 (
            .O(N__24758),
            .I(N__24749));
    InMux I__4861 (
            .O(N__24757),
            .I(N__24746));
    LocalMux I__4860 (
            .O(N__24754),
            .I(N__24743));
    Span4Mux_h I__4859 (
            .O(N__24749),
            .I(N__24740));
    LocalMux I__4858 (
            .O(N__24746),
            .I(N__24737));
    Sp12to4 I__4857 (
            .O(N__24743),
            .I(N__24734));
    Span4Mux_v I__4856 (
            .O(N__24740),
            .I(N__24731));
    Span4Mux_h I__4855 (
            .O(N__24737),
            .I(N__24726));
    Span12Mux_v I__4854 (
            .O(N__24734),
            .I(N__24723));
    Span4Mux_v I__4853 (
            .O(N__24731),
            .I(N__24720));
    InMux I__4852 (
            .O(N__24730),
            .I(N__24715));
    InMux I__4851 (
            .O(N__24729),
            .I(N__24715));
    Odrv4 I__4850 (
            .O(N__24726),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv12 I__4849 (
            .O(N__24723),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__4848 (
            .O(N__24720),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__4847 (
            .O(N__24715),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    InMux I__4846 (
            .O(N__24706),
            .I(N__24703));
    LocalMux I__4845 (
            .O(N__24703),
            .I(N__24695));
    InMux I__4844 (
            .O(N__24702),
            .I(N__24692));
    InMux I__4843 (
            .O(N__24701),
            .I(N__24689));
    InMux I__4842 (
            .O(N__24700),
            .I(N__24684));
    InMux I__4841 (
            .O(N__24699),
            .I(N__24684));
    InMux I__4840 (
            .O(N__24698),
            .I(N__24681));
    Span4Mux_v I__4839 (
            .O(N__24695),
            .I(N__24678));
    LocalMux I__4838 (
            .O(N__24692),
            .I(N__24675));
    LocalMux I__4837 (
            .O(N__24689),
            .I(N__24672));
    LocalMux I__4836 (
            .O(N__24684),
            .I(N__24669));
    LocalMux I__4835 (
            .O(N__24681),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__4834 (
            .O(N__24678),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv12 I__4833 (
            .O(N__24675),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__4832 (
            .O(N__24672),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv12 I__4831 (
            .O(N__24669),
            .I(M_this_oam_address_qZ0Z_1));
    InMux I__4830 (
            .O(N__24658),
            .I(N__24652));
    InMux I__4829 (
            .O(N__24657),
            .I(N__24649));
    InMux I__4828 (
            .O(N__24656),
            .I(N__24646));
    InMux I__4827 (
            .O(N__24655),
            .I(N__24640));
    LocalMux I__4826 (
            .O(N__24652),
            .I(N__24635));
    LocalMux I__4825 (
            .O(N__24649),
            .I(N__24635));
    LocalMux I__4824 (
            .O(N__24646),
            .I(N__24632));
    InMux I__4823 (
            .O(N__24645),
            .I(N__24627));
    InMux I__4822 (
            .O(N__24644),
            .I(N__24627));
    InMux I__4821 (
            .O(N__24643),
            .I(N__24624));
    LocalMux I__4820 (
            .O(N__24640),
            .I(N__24619));
    Span4Mux_v I__4819 (
            .O(N__24635),
            .I(N__24619));
    Span4Mux_v I__4818 (
            .O(N__24632),
            .I(N__24614));
    LocalMux I__4817 (
            .O(N__24627),
            .I(N__24614));
    LocalMux I__4816 (
            .O(N__24624),
            .I(N__24607));
    Span4Mux_v I__4815 (
            .O(N__24619),
            .I(N__24607));
    Span4Mux_v I__4814 (
            .O(N__24614),
            .I(N__24607));
    Odrv4 I__4813 (
            .O(N__24607),
            .I(M_this_oam_address_qZ0Z_0));
    CascadeMux I__4812 (
            .O(N__24604),
            .I(N__24599));
    CascadeMux I__4811 (
            .O(N__24603),
            .I(N__24596));
    InMux I__4810 (
            .O(N__24602),
            .I(N__24592));
    InMux I__4809 (
            .O(N__24599),
            .I(N__24589));
    InMux I__4808 (
            .O(N__24596),
            .I(N__24586));
    CascadeMux I__4807 (
            .O(N__24595),
            .I(N__24583));
    LocalMux I__4806 (
            .O(N__24592),
            .I(N__24575));
    LocalMux I__4805 (
            .O(N__24589),
            .I(N__24575));
    LocalMux I__4804 (
            .O(N__24586),
            .I(N__24575));
    InMux I__4803 (
            .O(N__24583),
            .I(N__24572));
    InMux I__4802 (
            .O(N__24582),
            .I(N__24568));
    Span4Mux_v I__4801 (
            .O(N__24575),
            .I(N__24565));
    LocalMux I__4800 (
            .O(N__24572),
            .I(N__24562));
    InMux I__4799 (
            .O(N__24571),
            .I(N__24559));
    LocalMux I__4798 (
            .O(N__24568),
            .I(N__24556));
    Span4Mux_h I__4797 (
            .O(N__24565),
            .I(N__24553));
    Sp12to4 I__4796 (
            .O(N__24562),
            .I(N__24548));
    LocalMux I__4795 (
            .O(N__24559),
            .I(N__24548));
    Odrv12 I__4794 (
            .O(N__24556),
            .I(N_314_1));
    Odrv4 I__4793 (
            .O(N__24553),
            .I(N_314_1));
    Odrv12 I__4792 (
            .O(N__24548),
            .I(N_314_1));
    CascadeMux I__4791 (
            .O(N__24541),
            .I(N__24537));
    InMux I__4790 (
            .O(N__24540),
            .I(N__24532));
    InMux I__4789 (
            .O(N__24537),
            .I(N__24532));
    LocalMux I__4788 (
            .O(N__24532),
            .I(N__24527));
    InMux I__4787 (
            .O(N__24531),
            .I(N__24524));
    InMux I__4786 (
            .O(N__24530),
            .I(N__24521));
    Span4Mux_v I__4785 (
            .O(N__24527),
            .I(N__24518));
    LocalMux I__4784 (
            .O(N__24524),
            .I(N__24515));
    LocalMux I__4783 (
            .O(N__24521),
            .I(N__24512));
    Span4Mux_h I__4782 (
            .O(N__24518),
            .I(N__24508));
    Span4Mux_v I__4781 (
            .O(N__24515),
            .I(N__24503));
    Span4Mux_v I__4780 (
            .O(N__24512),
            .I(N__24503));
    InMux I__4779 (
            .O(N__24511),
            .I(N__24500));
    Sp12to4 I__4778 (
            .O(N__24508),
            .I(N__24493));
    Sp12to4 I__4777 (
            .O(N__24503),
            .I(N__24493));
    LocalMux I__4776 (
            .O(N__24500),
            .I(N__24493));
    Span12Mux_h I__4775 (
            .O(N__24493),
            .I(N__24490));
    Odrv12 I__4774 (
            .O(N__24490),
            .I(port_enb_c));
    CascadeMux I__4773 (
            .O(N__24487),
            .I(N__24484));
    InMux I__4772 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__4771 (
            .O(N__24481),
            .I(N__24478));
    Span4Mux_v I__4770 (
            .O(N__24478),
            .I(N__24471));
    InMux I__4769 (
            .O(N__24477),
            .I(N__24468));
    InMux I__4768 (
            .O(N__24476),
            .I(N__24461));
    InMux I__4767 (
            .O(N__24475),
            .I(N__24461));
    InMux I__4766 (
            .O(N__24474),
            .I(N__24461));
    Odrv4 I__4765 (
            .O(N__24471),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__4764 (
            .O(N__24468),
            .I(this_start_data_delay_M_last_q));
    LocalMux I__4763 (
            .O(N__24461),
            .I(this_start_data_delay_M_last_q));
    InMux I__4762 (
            .O(N__24454),
            .I(N__24451));
    LocalMux I__4761 (
            .O(N__24451),
            .I(N__24446));
    InMux I__4760 (
            .O(N__24450),
            .I(N__24443));
    InMux I__4759 (
            .O(N__24449),
            .I(N__24438));
    Span4Mux_v I__4758 (
            .O(N__24446),
            .I(N__24433));
    LocalMux I__4757 (
            .O(N__24443),
            .I(N__24433));
    InMux I__4756 (
            .O(N__24442),
            .I(N__24428));
    InMux I__4755 (
            .O(N__24441),
            .I(N__24428));
    LocalMux I__4754 (
            .O(N__24438),
            .I(M_this_delay_clk_out_0));
    Odrv4 I__4753 (
            .O(N__24433),
            .I(M_this_delay_clk_out_0));
    LocalMux I__4752 (
            .O(N__24428),
            .I(M_this_delay_clk_out_0));
    CascadeMux I__4751 (
            .O(N__24421),
            .I(N_309_0_cascade_));
    InMux I__4750 (
            .O(N__24418),
            .I(N__24415));
    LocalMux I__4749 (
            .O(N__24415),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    InMux I__4748 (
            .O(N__24412),
            .I(N__24407));
    InMux I__4747 (
            .O(N__24411),
            .I(N__24404));
    InMux I__4746 (
            .O(N__24410),
            .I(N__24401));
    LocalMux I__4745 (
            .O(N__24407),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__4744 (
            .O(N__24404),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__4743 (
            .O(N__24401),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__4742 (
            .O(N__24394),
            .I(N__24391));
    LocalMux I__4741 (
            .O(N__24391),
            .I(M_this_data_count_q_cry_5_THRU_CO));
    CascadeMux I__4740 (
            .O(N__24388),
            .I(N__24383));
    InMux I__4739 (
            .O(N__24387),
            .I(N__24380));
    InMux I__4738 (
            .O(N__24386),
            .I(N__24377));
    InMux I__4737 (
            .O(N__24383),
            .I(N__24374));
    LocalMux I__4736 (
            .O(N__24380),
            .I(N__24371));
    LocalMux I__4735 (
            .O(N__24377),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__4734 (
            .O(N__24374),
            .I(M_this_data_count_qZ0Z_6));
    Odrv4 I__4733 (
            .O(N__24371),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__4732 (
            .O(N__24364),
            .I(N__24361));
    LocalMux I__4731 (
            .O(N__24361),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    CascadeMux I__4730 (
            .O(N__24358),
            .I(N__24353));
    CascadeMux I__4729 (
            .O(N__24357),
            .I(N__24350));
    InMux I__4728 (
            .O(N__24356),
            .I(N__24347));
    InMux I__4727 (
            .O(N__24353),
            .I(N__24344));
    InMux I__4726 (
            .O(N__24350),
            .I(N__24341));
    LocalMux I__4725 (
            .O(N__24347),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__4724 (
            .O(N__24344),
            .I(M_this_data_count_qZ0Z_7));
    LocalMux I__4723 (
            .O(N__24341),
            .I(M_this_data_count_qZ0Z_7));
    CascadeMux I__4722 (
            .O(N__24334),
            .I(N__24331));
    CascadeBuf I__4721 (
            .O(N__24331),
            .I(N__24328));
    CascadeMux I__4720 (
            .O(N__24328),
            .I(N__24325));
    InMux I__4719 (
            .O(N__24325),
            .I(N__24322));
    LocalMux I__4718 (
            .O(N__24322),
            .I(N__24319));
    Sp12to4 I__4717 (
            .O(N__24319),
            .I(N__24314));
    InMux I__4716 (
            .O(N__24318),
            .I(N__24311));
    InMux I__4715 (
            .O(N__24317),
            .I(N__24308));
    Span12Mux_h I__4714 (
            .O(N__24314),
            .I(N__24305));
    LocalMux I__4713 (
            .O(N__24311),
            .I(M_this_oam_address_qZ0Z_6));
    LocalMux I__4712 (
            .O(N__24308),
            .I(M_this_oam_address_qZ0Z_6));
    Odrv12 I__4711 (
            .O(N__24305),
            .I(M_this_oam_address_qZ0Z_6));
    CascadeMux I__4710 (
            .O(N__24298),
            .I(N__24295));
    CascadeBuf I__4709 (
            .O(N__24295),
            .I(N__24292));
    CascadeMux I__4708 (
            .O(N__24292),
            .I(N__24289));
    InMux I__4707 (
            .O(N__24289),
            .I(N__24286));
    LocalMux I__4706 (
            .O(N__24286),
            .I(N__24282));
    CascadeMux I__4705 (
            .O(N__24285),
            .I(N__24279));
    Span4Mux_h I__4704 (
            .O(N__24282),
            .I(N__24276));
    InMux I__4703 (
            .O(N__24279),
            .I(N__24273));
    Span4Mux_h I__4702 (
            .O(N__24276),
            .I(N__24270));
    LocalMux I__4701 (
            .O(N__24273),
            .I(N__24265));
    Span4Mux_v I__4700 (
            .O(N__24270),
            .I(N__24265));
    Odrv4 I__4699 (
            .O(N__24265),
            .I(M_this_oam_address_qZ0Z_7));
    InMux I__4698 (
            .O(N__24262),
            .I(N__24252));
    InMux I__4697 (
            .O(N__24261),
            .I(N__24249));
    InMux I__4696 (
            .O(N__24260),
            .I(N__24244));
    InMux I__4695 (
            .O(N__24259),
            .I(N__24244));
    InMux I__4694 (
            .O(N__24258),
            .I(N__24235));
    InMux I__4693 (
            .O(N__24257),
            .I(N__24235));
    InMux I__4692 (
            .O(N__24256),
            .I(N__24235));
    InMux I__4691 (
            .O(N__24255),
            .I(N__24235));
    LocalMux I__4690 (
            .O(N__24252),
            .I(N__24230));
    LocalMux I__4689 (
            .O(N__24249),
            .I(N__24223));
    LocalMux I__4688 (
            .O(N__24244),
            .I(N__24223));
    LocalMux I__4687 (
            .O(N__24235),
            .I(N__24223));
    InMux I__4686 (
            .O(N__24234),
            .I(N__24218));
    InMux I__4685 (
            .O(N__24233),
            .I(N__24218));
    Span4Mux_v I__4684 (
            .O(N__24230),
            .I(N__24215));
    Span4Mux_v I__4683 (
            .O(N__24223),
            .I(N__24210));
    LocalMux I__4682 (
            .O(N__24218),
            .I(N__24210));
    Sp12to4 I__4681 (
            .O(N__24215),
            .I(N__24207));
    Span4Mux_v I__4680 (
            .O(N__24210),
            .I(N__24204));
    Span12Mux_h I__4679 (
            .O(N__24207),
            .I(N__24201));
    Span4Mux_v I__4678 (
            .O(N__24204),
            .I(N__24198));
    Odrv12 I__4677 (
            .O(N__24201),
            .I(rst_n_c));
    Odrv4 I__4676 (
            .O(N__24198),
            .I(rst_n_c));
    InMux I__4675 (
            .O(N__24193),
            .I(N__24190));
    LocalMux I__4674 (
            .O(N__24190),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    InMux I__4673 (
            .O(N__24187),
            .I(N__24184));
    LocalMux I__4672 (
            .O(N__24184),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    CascadeMux I__4671 (
            .O(N__24181),
            .I(\this_ppu.N_760_0_cascade_ ));
    InMux I__4670 (
            .O(N__24178),
            .I(N__24175));
    LocalMux I__4669 (
            .O(N__24175),
            .I(N__24168));
    InMux I__4668 (
            .O(N__24174),
            .I(N__24165));
    InMux I__4667 (
            .O(N__24173),
            .I(N__24158));
    InMux I__4666 (
            .O(N__24172),
            .I(N__24158));
    InMux I__4665 (
            .O(N__24171),
            .I(N__24158));
    Span4Mux_v I__4664 (
            .O(N__24168),
            .I(N__24155));
    LocalMux I__4663 (
            .O(N__24165),
            .I(N__24150));
    LocalMux I__4662 (
            .O(N__24158),
            .I(N__24150));
    Span4Mux_v I__4661 (
            .O(N__24155),
            .I(N__24147));
    Span12Mux_h I__4660 (
            .O(N__24150),
            .I(N__24144));
    Span4Mux_h I__4659 (
            .O(N__24147),
            .I(N__24141));
    Span12Mux_v I__4658 (
            .O(N__24144),
            .I(N__24138));
    Odrv4 I__4657 (
            .O(N__24141),
            .I(\this_ppu.N_762_0 ));
    Odrv12 I__4656 (
            .O(N__24138),
            .I(\this_ppu.N_762_0 ));
    InMux I__4655 (
            .O(N__24133),
            .I(N__24130));
    LocalMux I__4654 (
            .O(N__24130),
            .I(N__24127));
    Span4Mux_h I__4653 (
            .O(N__24127),
            .I(N__24121));
    InMux I__4652 (
            .O(N__24126),
            .I(N__24118));
    InMux I__4651 (
            .O(N__24125),
            .I(N__24115));
    InMux I__4650 (
            .O(N__24124),
            .I(N__24112));
    Odrv4 I__4649 (
            .O(N__24121),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__4648 (
            .O(N__24118),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__4647 (
            .O(N__24115),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__4646 (
            .O(N__24112),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__4645 (
            .O(N__24103),
            .I(N__24100));
    InMux I__4644 (
            .O(N__24100),
            .I(N__24095));
    CascadeMux I__4643 (
            .O(N__24099),
            .I(N__24092));
    InMux I__4642 (
            .O(N__24098),
            .I(N__24089));
    LocalMux I__4641 (
            .O(N__24095),
            .I(N__24086));
    InMux I__4640 (
            .O(N__24092),
            .I(N__24082));
    LocalMux I__4639 (
            .O(N__24089),
            .I(N__24079));
    Span4Mux_v I__4638 (
            .O(N__24086),
            .I(N__24076));
    InMux I__4637 (
            .O(N__24085),
            .I(N__24073));
    LocalMux I__4636 (
            .O(N__24082),
            .I(N__24070));
    Sp12to4 I__4635 (
            .O(N__24079),
            .I(N__24067));
    Span4Mux_v I__4634 (
            .O(N__24076),
            .I(N__24063));
    LocalMux I__4633 (
            .O(N__24073),
            .I(N__24058));
    Span4Mux_h I__4632 (
            .O(N__24070),
            .I(N__24058));
    Span12Mux_v I__4631 (
            .O(N__24067),
            .I(N__24055));
    InMux I__4630 (
            .O(N__24066),
            .I(N__24052));
    Odrv4 I__4629 (
            .O(N__24063),
            .I(\this_ppu.M_last_q ));
    Odrv4 I__4628 (
            .O(N__24058),
            .I(\this_ppu.M_last_q ));
    Odrv12 I__4627 (
            .O(N__24055),
            .I(\this_ppu.M_last_q ));
    LocalMux I__4626 (
            .O(N__24052),
            .I(\this_ppu.M_last_q ));
    InMux I__4625 (
            .O(N__24043),
            .I(N__24040));
    LocalMux I__4624 (
            .O(N__24040),
            .I(N__24035));
    InMux I__4623 (
            .O(N__24039),
            .I(N__24032));
    InMux I__4622 (
            .O(N__24038),
            .I(N__24028));
    Span4Mux_h I__4621 (
            .O(N__24035),
            .I(N__24023));
    LocalMux I__4620 (
            .O(N__24032),
            .I(N__24023));
    InMux I__4619 (
            .O(N__24031),
            .I(N__24020));
    LocalMux I__4618 (
            .O(N__24028),
            .I(N__24017));
    Span4Mux_v I__4617 (
            .O(N__24023),
            .I(N__24014));
    LocalMux I__4616 (
            .O(N__24020),
            .I(N__24009));
    Span4Mux_h I__4615 (
            .O(N__24017),
            .I(N__24009));
    Span4Mux_h I__4614 (
            .O(N__24014),
            .I(N__24006));
    Odrv4 I__4613 (
            .O(N__24009),
            .I(\this_ppu.N_5_4 ));
    Odrv4 I__4612 (
            .O(N__24006),
            .I(\this_ppu.N_5_4 ));
    InMux I__4611 (
            .O(N__24001),
            .I(N__23998));
    LocalMux I__4610 (
            .O(N__23998),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ));
    CascadeMux I__4609 (
            .O(N__23995),
            .I(\this_ppu.N_268_i_0_0_cascade_ ));
    InMux I__4608 (
            .O(N__23992),
            .I(N__23987));
    InMux I__4607 (
            .O(N__23991),
            .I(N__23984));
    InMux I__4606 (
            .O(N__23990),
            .I(N__23981));
    LocalMux I__4605 (
            .O(N__23987),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__4604 (
            .O(N__23984),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    LocalMux I__4603 (
            .O(N__23981),
            .I(\this_ppu.M_count_qZ0Z_5 ));
    IoInMux I__4602 (
            .O(N__23974),
            .I(N__23970));
    InMux I__4601 (
            .O(N__23973),
            .I(N__23967));
    LocalMux I__4600 (
            .O(N__23970),
            .I(N__23964));
    LocalMux I__4599 (
            .O(N__23967),
            .I(N__23961));
    IoSpan4Mux I__4598 (
            .O(N__23964),
            .I(N__23950));
    Span4Mux_v I__4597 (
            .O(N__23961),
            .I(N__23947));
    InMux I__4596 (
            .O(N__23960),
            .I(N__23938));
    InMux I__4595 (
            .O(N__23959),
            .I(N__23938));
    InMux I__4594 (
            .O(N__23958),
            .I(N__23938));
    InMux I__4593 (
            .O(N__23957),
            .I(N__23938));
    InMux I__4592 (
            .O(N__23956),
            .I(N__23933));
    InMux I__4591 (
            .O(N__23955),
            .I(N__23933));
    InMux I__4590 (
            .O(N__23954),
            .I(N__23930));
    InMux I__4589 (
            .O(N__23953),
            .I(N__23927));
    Span4Mux_s1_h I__4588 (
            .O(N__23950),
            .I(N__23924));
    Sp12to4 I__4587 (
            .O(N__23947),
            .I(N__23919));
    LocalMux I__4586 (
            .O(N__23938),
            .I(N__23919));
    LocalMux I__4585 (
            .O(N__23933),
            .I(N__23916));
    LocalMux I__4584 (
            .O(N__23930),
            .I(N__23913));
    LocalMux I__4583 (
            .O(N__23927),
            .I(N__23910));
    Sp12to4 I__4582 (
            .O(N__23924),
            .I(N__23907));
    Span12Mux_h I__4581 (
            .O(N__23919),
            .I(N__23904));
    Span12Mux_s11_h I__4580 (
            .O(N__23916),
            .I(N__23899));
    Span12Mux_v I__4579 (
            .O(N__23913),
            .I(N__23899));
    Span12Mux_v I__4578 (
            .O(N__23910),
            .I(N__23894));
    Span12Mux_h I__4577 (
            .O(N__23907),
            .I(N__23894));
    Odrv12 I__4576 (
            .O(N__23904),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__4575 (
            .O(N__23899),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__4574 (
            .O(N__23894),
            .I(M_this_reset_cond_out_0));
    InMux I__4573 (
            .O(N__23887),
            .I(N__23884));
    LocalMux I__4572 (
            .O(N__23884),
            .I(N__23881));
    Odrv4 I__4571 (
            .O(N__23881),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ));
    CascadeMux I__4570 (
            .O(N__23878),
            .I(\this_ppu.N_1323_0_cascade_ ));
    InMux I__4569 (
            .O(N__23875),
            .I(N__23870));
    InMux I__4568 (
            .O(N__23874),
            .I(N__23867));
    InMux I__4567 (
            .O(N__23873),
            .I(N__23864));
    LocalMux I__4566 (
            .O(N__23870),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__4565 (
            .O(N__23867),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    LocalMux I__4564 (
            .O(N__23864),
            .I(\this_ppu.M_count_qZ0Z_1 ));
    InMux I__4563 (
            .O(N__23857),
            .I(N__23853));
    InMux I__4562 (
            .O(N__23856),
            .I(N__23850));
    LocalMux I__4561 (
            .O(N__23853),
            .I(N__23845));
    LocalMux I__4560 (
            .O(N__23850),
            .I(N__23845));
    Odrv4 I__4559 (
            .O(N__23845),
            .I(\this_ppu.M_count_qZ0Z_7 ));
    InMux I__4558 (
            .O(N__23842),
            .I(N__23839));
    LocalMux I__4557 (
            .O(N__23839),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3 ));
    InMux I__4556 (
            .O(N__23836),
            .I(bfn_17_19_0_));
    InMux I__4555 (
            .O(N__23833),
            .I(N__23830));
    LocalMux I__4554 (
            .O(N__23830),
            .I(N__23827));
    Odrv4 I__4553 (
            .O(N__23827),
            .I(M_this_data_count_q_cry_8_THRU_CO));
    InMux I__4552 (
            .O(N__23824),
            .I(M_this_data_count_q_cry_8));
    InMux I__4551 (
            .O(N__23821),
            .I(N__23817));
    InMux I__4550 (
            .O(N__23820),
            .I(N__23814));
    LocalMux I__4549 (
            .O(N__23817),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__4548 (
            .O(N__23814),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__4547 (
            .O(N__23809),
            .I(N__23806));
    LocalMux I__4546 (
            .O(N__23806),
            .I(M_this_data_count_q_s_10));
    InMux I__4545 (
            .O(N__23803),
            .I(M_this_data_count_q_cry_9));
    CascadeMux I__4544 (
            .O(N__23800),
            .I(N__23797));
    InMux I__4543 (
            .O(N__23797),
            .I(N__23792));
    InMux I__4542 (
            .O(N__23796),
            .I(N__23787));
    InMux I__4541 (
            .O(N__23795),
            .I(N__23787));
    LocalMux I__4540 (
            .O(N__23792),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__4539 (
            .O(N__23787),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__4538 (
            .O(N__23782),
            .I(N__23779));
    InMux I__4537 (
            .O(N__23779),
            .I(N__23776));
    LocalMux I__4536 (
            .O(N__23776),
            .I(M_this_data_count_q_cry_10_THRU_CO));
    InMux I__4535 (
            .O(N__23773),
            .I(M_this_data_count_q_cry_10));
    CascadeMux I__4534 (
            .O(N__23770),
            .I(N__23764));
    CascadeMux I__4533 (
            .O(N__23769),
            .I(N__23760));
    CascadeMux I__4532 (
            .O(N__23768),
            .I(N__23756));
    InMux I__4531 (
            .O(N__23767),
            .I(N__23736));
    InMux I__4530 (
            .O(N__23764),
            .I(N__23736));
    InMux I__4529 (
            .O(N__23763),
            .I(N__23736));
    InMux I__4528 (
            .O(N__23760),
            .I(N__23736));
    InMux I__4527 (
            .O(N__23759),
            .I(N__23736));
    InMux I__4526 (
            .O(N__23756),
            .I(N__23736));
    CascadeMux I__4525 (
            .O(N__23755),
            .I(N__23732));
    CascadeMux I__4524 (
            .O(N__23754),
            .I(N__23729));
    SRMux I__4523 (
            .O(N__23753),
            .I(N__23726));
    SRMux I__4522 (
            .O(N__23752),
            .I(N__23723));
    SRMux I__4521 (
            .O(N__23751),
            .I(N__23720));
    IoInMux I__4520 (
            .O(N__23750),
            .I(N__23714));
    CascadeMux I__4519 (
            .O(N__23749),
            .I(N__23709));
    LocalMux I__4518 (
            .O(N__23736),
            .I(N__23705));
    InMux I__4517 (
            .O(N__23735),
            .I(N__23698));
    InMux I__4516 (
            .O(N__23732),
            .I(N__23698));
    InMux I__4515 (
            .O(N__23729),
            .I(N__23698));
    LocalMux I__4514 (
            .O(N__23726),
            .I(N__23689));
    LocalMux I__4513 (
            .O(N__23723),
            .I(N__23689));
    LocalMux I__4512 (
            .O(N__23720),
            .I(N__23686));
    SRMux I__4511 (
            .O(N__23719),
            .I(N__23683));
    SRMux I__4510 (
            .O(N__23718),
            .I(N__23680));
    SRMux I__4509 (
            .O(N__23717),
            .I(N__23677));
    LocalMux I__4508 (
            .O(N__23714),
            .I(N__23671));
    SRMux I__4507 (
            .O(N__23713),
            .I(N__23668));
    SRMux I__4506 (
            .O(N__23712),
            .I(N__23664));
    InMux I__4505 (
            .O(N__23709),
            .I(N__23657));
    InMux I__4504 (
            .O(N__23708),
            .I(N__23657));
    Span4Mux_h I__4503 (
            .O(N__23705),
            .I(N__23652));
    LocalMux I__4502 (
            .O(N__23698),
            .I(N__23652));
    InMux I__4501 (
            .O(N__23697),
            .I(N__23649));
    CascadeMux I__4500 (
            .O(N__23696),
            .I(N__23645));
    CascadeMux I__4499 (
            .O(N__23695),
            .I(N__23641));
    CascadeMux I__4498 (
            .O(N__23694),
            .I(N__23637));
    Span4Mux_v I__4497 (
            .O(N__23689),
            .I(N__23627));
    Span4Mux_h I__4496 (
            .O(N__23686),
            .I(N__23627));
    LocalMux I__4495 (
            .O(N__23683),
            .I(N__23627));
    LocalMux I__4494 (
            .O(N__23680),
            .I(N__23627));
    LocalMux I__4493 (
            .O(N__23677),
            .I(N__23624));
    SRMux I__4492 (
            .O(N__23676),
            .I(N__23621));
    SRMux I__4491 (
            .O(N__23675),
            .I(N__23618));
    SRMux I__4490 (
            .O(N__23674),
            .I(N__23615));
    IoSpan4Mux I__4489 (
            .O(N__23671),
            .I(N__23610));
    LocalMux I__4488 (
            .O(N__23668),
            .I(N__23607));
    SRMux I__4487 (
            .O(N__23667),
            .I(N__23604));
    LocalMux I__4486 (
            .O(N__23664),
            .I(N__23601));
    SRMux I__4485 (
            .O(N__23663),
            .I(N__23598));
    SRMux I__4484 (
            .O(N__23662),
            .I(N__23592));
    LocalMux I__4483 (
            .O(N__23657),
            .I(N__23588));
    Span4Mux_v I__4482 (
            .O(N__23652),
            .I(N__23583));
    LocalMux I__4481 (
            .O(N__23649),
            .I(N__23583));
    InMux I__4480 (
            .O(N__23648),
            .I(N__23570));
    InMux I__4479 (
            .O(N__23645),
            .I(N__23570));
    InMux I__4478 (
            .O(N__23644),
            .I(N__23570));
    InMux I__4477 (
            .O(N__23641),
            .I(N__23570));
    InMux I__4476 (
            .O(N__23640),
            .I(N__23570));
    InMux I__4475 (
            .O(N__23637),
            .I(N__23570));
    IoInMux I__4474 (
            .O(N__23636),
            .I(N__23567));
    Span4Mux_v I__4473 (
            .O(N__23627),
            .I(N__23558));
    Span4Mux_h I__4472 (
            .O(N__23624),
            .I(N__23558));
    LocalMux I__4471 (
            .O(N__23621),
            .I(N__23558));
    LocalMux I__4470 (
            .O(N__23618),
            .I(N__23558));
    LocalMux I__4469 (
            .O(N__23615),
            .I(N__23555));
    SRMux I__4468 (
            .O(N__23614),
            .I(N__23552));
    SRMux I__4467 (
            .O(N__23613),
            .I(N__23549));
    Span4Mux_s3_h I__4466 (
            .O(N__23610),
            .I(N__23542));
    Span4Mux_v I__4465 (
            .O(N__23607),
            .I(N__23537));
    LocalMux I__4464 (
            .O(N__23604),
            .I(N__23537));
    Span4Mux_v I__4463 (
            .O(N__23601),
            .I(N__23532));
    LocalMux I__4462 (
            .O(N__23598),
            .I(N__23532));
    SRMux I__4461 (
            .O(N__23597),
            .I(N__23529));
    SRMux I__4460 (
            .O(N__23596),
            .I(N__23526));
    SRMux I__4459 (
            .O(N__23595),
            .I(N__23518));
    LocalMux I__4458 (
            .O(N__23592),
            .I(N__23515));
    SRMux I__4457 (
            .O(N__23591),
            .I(N__23510));
    Span4Mux_v I__4456 (
            .O(N__23588),
            .I(N__23503));
    Span4Mux_h I__4455 (
            .O(N__23583),
            .I(N__23503));
    LocalMux I__4454 (
            .O(N__23570),
            .I(N__23503));
    LocalMux I__4453 (
            .O(N__23567),
            .I(N__23500));
    Span4Mux_v I__4452 (
            .O(N__23558),
            .I(N__23491));
    Span4Mux_h I__4451 (
            .O(N__23555),
            .I(N__23491));
    LocalMux I__4450 (
            .O(N__23552),
            .I(N__23491));
    LocalMux I__4449 (
            .O(N__23549),
            .I(N__23491));
    SRMux I__4448 (
            .O(N__23548),
            .I(N__23488));
    SRMux I__4447 (
            .O(N__23547),
            .I(N__23485));
    SRMux I__4446 (
            .O(N__23546),
            .I(N__23482));
    SRMux I__4445 (
            .O(N__23545),
            .I(N__23478));
    Span4Mux_h I__4444 (
            .O(N__23542),
            .I(N__23466));
    Span4Mux_v I__4443 (
            .O(N__23537),
            .I(N__23466));
    Span4Mux_v I__4442 (
            .O(N__23532),
            .I(N__23466));
    LocalMux I__4441 (
            .O(N__23529),
            .I(N__23466));
    LocalMux I__4440 (
            .O(N__23526),
            .I(N__23463));
    SRMux I__4439 (
            .O(N__23525),
            .I(N__23460));
    SRMux I__4438 (
            .O(N__23524),
            .I(N__23457));
    SRMux I__4437 (
            .O(N__23523),
            .I(N__23451));
    SRMux I__4436 (
            .O(N__23522),
            .I(N__23448));
    SRMux I__4435 (
            .O(N__23521),
            .I(N__23442));
    LocalMux I__4434 (
            .O(N__23518),
            .I(N__23437));
    Span4Mux_h I__4433 (
            .O(N__23515),
            .I(N__23437));
    SRMux I__4432 (
            .O(N__23514),
            .I(N__23434));
    SRMux I__4431 (
            .O(N__23513),
            .I(N__23431));
    LocalMux I__4430 (
            .O(N__23510),
            .I(N__23425));
    Span4Mux_v I__4429 (
            .O(N__23503),
            .I(N__23422));
    Span4Mux_s2_h I__4428 (
            .O(N__23500),
            .I(N__23419));
    Span4Mux_v I__4427 (
            .O(N__23491),
            .I(N__23412));
    LocalMux I__4426 (
            .O(N__23488),
            .I(N__23412));
    LocalMux I__4425 (
            .O(N__23485),
            .I(N__23412));
    LocalMux I__4424 (
            .O(N__23482),
            .I(N__23409));
    SRMux I__4423 (
            .O(N__23481),
            .I(N__23406));
    LocalMux I__4422 (
            .O(N__23478),
            .I(N__23402));
    SRMux I__4421 (
            .O(N__23477),
            .I(N__23399));
    SRMux I__4420 (
            .O(N__23476),
            .I(N__23396));
    SRMux I__4419 (
            .O(N__23475),
            .I(N__23393));
    Span4Mux_v I__4418 (
            .O(N__23466),
            .I(N__23384));
    Span4Mux_v I__4417 (
            .O(N__23463),
            .I(N__23384));
    LocalMux I__4416 (
            .O(N__23460),
            .I(N__23384));
    LocalMux I__4415 (
            .O(N__23457),
            .I(N__23384));
    SRMux I__4414 (
            .O(N__23456),
            .I(N__23381));
    SRMux I__4413 (
            .O(N__23455),
            .I(N__23378));
    SRMux I__4412 (
            .O(N__23454),
            .I(N__23375));
    LocalMux I__4411 (
            .O(N__23451),
            .I(N__23370));
    LocalMux I__4410 (
            .O(N__23448),
            .I(N__23370));
    SRMux I__4409 (
            .O(N__23447),
            .I(N__23367));
    SRMux I__4408 (
            .O(N__23446),
            .I(N__23364));
    SRMux I__4407 (
            .O(N__23445),
            .I(N__23360));
    LocalMux I__4406 (
            .O(N__23442),
            .I(N__23351));
    Sp12to4 I__4405 (
            .O(N__23437),
            .I(N__23351));
    LocalMux I__4404 (
            .O(N__23434),
            .I(N__23351));
    LocalMux I__4403 (
            .O(N__23431),
            .I(N__23351));
    SRMux I__4402 (
            .O(N__23430),
            .I(N__23348));
    SRMux I__4401 (
            .O(N__23429),
            .I(N__23345));
    SRMux I__4400 (
            .O(N__23428),
            .I(N__23342));
    Span4Mux_h I__4399 (
            .O(N__23425),
            .I(N__23339));
    Span4Mux_v I__4398 (
            .O(N__23422),
            .I(N__23336));
    Span4Mux_h I__4397 (
            .O(N__23419),
            .I(N__23331));
    Span4Mux_v I__4396 (
            .O(N__23412),
            .I(N__23331));
    Span4Mux_h I__4395 (
            .O(N__23409),
            .I(N__23328));
    LocalMux I__4394 (
            .O(N__23406),
            .I(N__23325));
    SRMux I__4393 (
            .O(N__23405),
            .I(N__23322));
    Span4Mux_s1_v I__4392 (
            .O(N__23402),
            .I(N__23315));
    LocalMux I__4391 (
            .O(N__23399),
            .I(N__23315));
    LocalMux I__4390 (
            .O(N__23396),
            .I(N__23315));
    LocalMux I__4389 (
            .O(N__23393),
            .I(N__23312));
    Span4Mux_v I__4388 (
            .O(N__23384),
            .I(N__23305));
    LocalMux I__4387 (
            .O(N__23381),
            .I(N__23305));
    LocalMux I__4386 (
            .O(N__23378),
            .I(N__23305));
    LocalMux I__4385 (
            .O(N__23375),
            .I(N__23302));
    Span4Mux_v I__4384 (
            .O(N__23370),
            .I(N__23295));
    LocalMux I__4383 (
            .O(N__23367),
            .I(N__23295));
    LocalMux I__4382 (
            .O(N__23364),
            .I(N__23295));
    SRMux I__4381 (
            .O(N__23363),
            .I(N__23292));
    LocalMux I__4380 (
            .O(N__23360),
            .I(N__23289));
    Span12Mux_v I__4379 (
            .O(N__23351),
            .I(N__23280));
    LocalMux I__4378 (
            .O(N__23348),
            .I(N__23280));
    LocalMux I__4377 (
            .O(N__23345),
            .I(N__23280));
    LocalMux I__4376 (
            .O(N__23342),
            .I(N__23280));
    Span4Mux_v I__4375 (
            .O(N__23339),
            .I(N__23273));
    Span4Mux_v I__4374 (
            .O(N__23336),
            .I(N__23273));
    Span4Mux_h I__4373 (
            .O(N__23331),
            .I(N__23273));
    Span4Mux_v I__4372 (
            .O(N__23328),
            .I(N__23268));
    Span4Mux_h I__4371 (
            .O(N__23325),
            .I(N__23268));
    LocalMux I__4370 (
            .O(N__23322),
            .I(N__23263));
    Sp12to4 I__4369 (
            .O(N__23315),
            .I(N__23263));
    Span4Mux_v I__4368 (
            .O(N__23312),
            .I(N__23258));
    Span4Mux_v I__4367 (
            .O(N__23305),
            .I(N__23258));
    Span4Mux_v I__4366 (
            .O(N__23302),
            .I(N__23251));
    Span4Mux_v I__4365 (
            .O(N__23295),
            .I(N__23251));
    LocalMux I__4364 (
            .O(N__23292),
            .I(N__23251));
    Span4Mux_h I__4363 (
            .O(N__23289),
            .I(N__23248));
    Span12Mux_v I__4362 (
            .O(N__23280),
            .I(N__23239));
    Sp12to4 I__4361 (
            .O(N__23273),
            .I(N__23239));
    Sp12to4 I__4360 (
            .O(N__23268),
            .I(N__23239));
    Span12Mux_s5_v I__4359 (
            .O(N__23263),
            .I(N__23239));
    Span4Mux_h I__4358 (
            .O(N__23258),
            .I(N__23234));
    Span4Mux_h I__4357 (
            .O(N__23251),
            .I(N__23234));
    Span4Mux_h I__4356 (
            .O(N__23248),
            .I(N__23231));
    Odrv12 I__4355 (
            .O(N__23239),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4354 (
            .O(N__23234),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4353 (
            .O(N__23231),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__4352 (
            .O(N__23224),
            .I(N__23221));
    InMux I__4351 (
            .O(N__23221),
            .I(N__23216));
    InMux I__4350 (
            .O(N__23220),
            .I(N__23211));
    InMux I__4349 (
            .O(N__23219),
            .I(N__23211));
    LocalMux I__4348 (
            .O(N__23216),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__4347 (
            .O(N__23211),
            .I(M_this_data_count_qZ0Z_12));
    InMux I__4346 (
            .O(N__23206),
            .I(N__23203));
    LocalMux I__4345 (
            .O(N__23203),
            .I(M_this_data_count_q_cry_11_THRU_CO));
    InMux I__4344 (
            .O(N__23200),
            .I(M_this_data_count_q_cry_11));
    InMux I__4343 (
            .O(N__23197),
            .I(M_this_data_count_q_cry_12));
    InMux I__4342 (
            .O(N__23194),
            .I(N__23189));
    InMux I__4341 (
            .O(N__23193),
            .I(N__23186));
    InMux I__4340 (
            .O(N__23192),
            .I(N__23183));
    LocalMux I__4339 (
            .O(N__23189),
            .I(N__23180));
    LocalMux I__4338 (
            .O(N__23186),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__4337 (
            .O(N__23183),
            .I(M_this_data_count_qZ0Z_5));
    Odrv4 I__4336 (
            .O(N__23180),
            .I(M_this_data_count_qZ0Z_5));
    CascadeMux I__4335 (
            .O(N__23173),
            .I(N__23169));
    InMux I__4334 (
            .O(N__23172),
            .I(N__23163));
    InMux I__4333 (
            .O(N__23169),
            .I(N__23163));
    InMux I__4332 (
            .O(N__23168),
            .I(N__23160));
    LocalMux I__4331 (
            .O(N__23163),
            .I(N__23157));
    LocalMux I__4330 (
            .O(N__23160),
            .I(M_this_data_count_qZ0Z_9));
    Odrv4 I__4329 (
            .O(N__23157),
            .I(M_this_data_count_qZ0Z_9));
    CascadeMux I__4328 (
            .O(N__23152),
            .I(N__23149));
    InMux I__4327 (
            .O(N__23149),
            .I(N__23144));
    InMux I__4326 (
            .O(N__23148),
            .I(N__23141));
    InMux I__4325 (
            .O(N__23147),
            .I(N__23138));
    LocalMux I__4324 (
            .O(N__23144),
            .I(N__23133));
    LocalMux I__4323 (
            .O(N__23141),
            .I(N__23133));
    LocalMux I__4322 (
            .O(N__23138),
            .I(M_this_data_count_qZ0Z_4));
    Odrv4 I__4321 (
            .O(N__23133),
            .I(M_this_data_count_qZ0Z_4));
    InMux I__4320 (
            .O(N__23128),
            .I(N__23125));
    LocalMux I__4319 (
            .O(N__23125),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11 ));
    InMux I__4318 (
            .O(N__23122),
            .I(N__23119));
    LocalMux I__4317 (
            .O(N__23119),
            .I(N__23116));
    Span4Mux_h I__4316 (
            .O(N__23116),
            .I(N__23111));
    InMux I__4315 (
            .O(N__23115),
            .I(N__23106));
    InMux I__4314 (
            .O(N__23114),
            .I(N__23106));
    Odrv4 I__4313 (
            .O(N__23111),
            .I(\this_ppu.N_91 ));
    LocalMux I__4312 (
            .O(N__23106),
            .I(\this_ppu.N_91 ));
    InMux I__4311 (
            .O(N__23101),
            .I(N__23098));
    LocalMux I__4310 (
            .O(N__23098),
            .I(N__23095));
    Odrv4 I__4309 (
            .O(N__23095),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11 ));
    InMux I__4308 (
            .O(N__23092),
            .I(N__23087));
    InMux I__4307 (
            .O(N__23091),
            .I(N__23082));
    InMux I__4306 (
            .O(N__23090),
            .I(N__23082));
    LocalMux I__4305 (
            .O(N__23087),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__4304 (
            .O(N__23082),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__4303 (
            .O(N__23077),
            .I(M_this_data_count_q_cry_0));
    CascadeMux I__4302 (
            .O(N__23074),
            .I(N__23071));
    InMux I__4301 (
            .O(N__23071),
            .I(N__23066));
    InMux I__4300 (
            .O(N__23070),
            .I(N__23061));
    InMux I__4299 (
            .O(N__23069),
            .I(N__23061));
    LocalMux I__4298 (
            .O(N__23066),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__4297 (
            .O(N__23061),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__4296 (
            .O(N__23056),
            .I(N__23053));
    LocalMux I__4295 (
            .O(N__23053),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    InMux I__4294 (
            .O(N__23050),
            .I(M_this_data_count_q_cry_1));
    InMux I__4293 (
            .O(N__23047),
            .I(N__23042));
    InMux I__4292 (
            .O(N__23046),
            .I(N__23039));
    InMux I__4291 (
            .O(N__23045),
            .I(N__23036));
    LocalMux I__4290 (
            .O(N__23042),
            .I(N__23033));
    LocalMux I__4289 (
            .O(N__23039),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__4288 (
            .O(N__23036),
            .I(M_this_data_count_qZ0Z_3));
    Odrv4 I__4287 (
            .O(N__23033),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__4286 (
            .O(N__23026),
            .I(N__23023));
    LocalMux I__4285 (
            .O(N__23023),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    InMux I__4284 (
            .O(N__23020),
            .I(M_this_data_count_q_cry_2));
    InMux I__4283 (
            .O(N__23017),
            .I(N__23014));
    LocalMux I__4282 (
            .O(N__23014),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    InMux I__4281 (
            .O(N__23011),
            .I(M_this_data_count_q_cry_3));
    InMux I__4280 (
            .O(N__23008),
            .I(N__23005));
    LocalMux I__4279 (
            .O(N__23005),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    InMux I__4278 (
            .O(N__23002),
            .I(M_this_data_count_q_cry_4));
    InMux I__4277 (
            .O(N__22999),
            .I(M_this_data_count_q_cry_5));
    InMux I__4276 (
            .O(N__22996),
            .I(M_this_data_count_q_cry_6));
    InMux I__4275 (
            .O(N__22993),
            .I(N__22990));
    LocalMux I__4274 (
            .O(N__22990),
            .I(N__22987));
    Span4Mux_v I__4273 (
            .O(N__22987),
            .I(N__22984));
    Span4Mux_h I__4272 (
            .O(N__22984),
            .I(N__22981));
    Span4Mux_h I__4271 (
            .O(N__22981),
            .I(N__22978));
    Odrv4 I__4270 (
            .O(N__22978),
            .I(\this_ppu.oam_cache.mem_5 ));
    InMux I__4269 (
            .O(N__22975),
            .I(N__22972));
    LocalMux I__4268 (
            .O(N__22972),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_5 ));
    InMux I__4267 (
            .O(N__22969),
            .I(N__22965));
    InMux I__4266 (
            .O(N__22968),
            .I(N__22961));
    LocalMux I__4265 (
            .O(N__22965),
            .I(N__22957));
    InMux I__4264 (
            .O(N__22964),
            .I(N__22954));
    LocalMux I__4263 (
            .O(N__22961),
            .I(N__22950));
    InMux I__4262 (
            .O(N__22960),
            .I(N__22947));
    Span4Mux_h I__4261 (
            .O(N__22957),
            .I(N__22942));
    LocalMux I__4260 (
            .O(N__22954),
            .I(N__22939));
    InMux I__4259 (
            .O(N__22953),
            .I(N__22936));
    Span4Mux_h I__4258 (
            .O(N__22950),
            .I(N__22933));
    LocalMux I__4257 (
            .O(N__22947),
            .I(N__22930));
    InMux I__4256 (
            .O(N__22946),
            .I(N__22927));
    InMux I__4255 (
            .O(N__22945),
            .I(N__22923));
    Span4Mux_v I__4254 (
            .O(N__22942),
            .I(N__22918));
    Span4Mux_h I__4253 (
            .O(N__22939),
            .I(N__22918));
    LocalMux I__4252 (
            .O(N__22936),
            .I(N__22915));
    Span4Mux_v I__4251 (
            .O(N__22933),
            .I(N__22910));
    Span4Mux_h I__4250 (
            .O(N__22930),
            .I(N__22910));
    LocalMux I__4249 (
            .O(N__22927),
            .I(N__22907));
    InMux I__4248 (
            .O(N__22926),
            .I(N__22904));
    LocalMux I__4247 (
            .O(N__22923),
            .I(N__22901));
    Span4Mux_v I__4246 (
            .O(N__22918),
            .I(N__22896));
    Span4Mux_h I__4245 (
            .O(N__22915),
            .I(N__22896));
    Span4Mux_v I__4244 (
            .O(N__22910),
            .I(N__22891));
    Span4Mux_h I__4243 (
            .O(N__22907),
            .I(N__22891));
    LocalMux I__4242 (
            .O(N__22904),
            .I(N__22888));
    Span4Mux_h I__4241 (
            .O(N__22901),
            .I(N__22885));
    Span4Mux_h I__4240 (
            .O(N__22896),
            .I(N__22882));
    Span4Mux_v I__4239 (
            .O(N__22891),
            .I(N__22877));
    Span4Mux_h I__4238 (
            .O(N__22888),
            .I(N__22877));
    Span4Mux_h I__4237 (
            .O(N__22885),
            .I(N__22870));
    Span4Mux_h I__4236 (
            .O(N__22882),
            .I(N__22870));
    Span4Mux_h I__4235 (
            .O(N__22877),
            .I(N__22870));
    Odrv4 I__4234 (
            .O(N__22870),
            .I(M_this_spr_ram_write_data_1));
    InMux I__4233 (
            .O(N__22867),
            .I(N__22853));
    InMux I__4232 (
            .O(N__22866),
            .I(N__22853));
    InMux I__4231 (
            .O(N__22865),
            .I(N__22844));
    InMux I__4230 (
            .O(N__22864),
            .I(N__22844));
    InMux I__4229 (
            .O(N__22863),
            .I(N__22844));
    InMux I__4228 (
            .O(N__22862),
            .I(N__22844));
    InMux I__4227 (
            .O(N__22861),
            .I(N__22835));
    InMux I__4226 (
            .O(N__22860),
            .I(N__22835));
    InMux I__4225 (
            .O(N__22859),
            .I(N__22835));
    InMux I__4224 (
            .O(N__22858),
            .I(N__22835));
    LocalMux I__4223 (
            .O(N__22853),
            .I(N__22828));
    LocalMux I__4222 (
            .O(N__22844),
            .I(N__22828));
    LocalMux I__4221 (
            .O(N__22835),
            .I(N__22828));
    Span4Mux_v I__4220 (
            .O(N__22828),
            .I(N__22824));
    InMux I__4219 (
            .O(N__22827),
            .I(N__22821));
    Span4Mux_h I__4218 (
            .O(N__22824),
            .I(N__22818));
    LocalMux I__4217 (
            .O(N__22821),
            .I(N__22813));
    Span4Mux_h I__4216 (
            .O(N__22818),
            .I(N__22813));
    Odrv4 I__4215 (
            .O(N__22813),
            .I(N_609));
    InMux I__4214 (
            .O(N__22810),
            .I(N__22807));
    LocalMux I__4213 (
            .O(N__22807),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    InMux I__4212 (
            .O(N__22804),
            .I(N__22801));
    LocalMux I__4211 (
            .O(N__22801),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__4210 (
            .O(N__22798),
            .I(N__22795));
    LocalMux I__4209 (
            .O(N__22795),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__4208 (
            .O(N__22792),
            .I(N__22789));
    LocalMux I__4207 (
            .O(N__22789),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    InMux I__4206 (
            .O(N__22786),
            .I(N__22783));
    LocalMux I__4205 (
            .O(N__22783),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__4204 (
            .O(N__22780),
            .I(N__22777));
    LocalMux I__4203 (
            .O(N__22777),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__4202 (
            .O(N__22774),
            .I(N__22771));
    LocalMux I__4201 (
            .O(N__22771),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CEMux I__4200 (
            .O(N__22768),
            .I(N__22765));
    LocalMux I__4199 (
            .O(N__22765),
            .I(N__22761));
    CEMux I__4198 (
            .O(N__22764),
            .I(N__22758));
    Span4Mux_v I__4197 (
            .O(N__22761),
            .I(N__22753));
    LocalMux I__4196 (
            .O(N__22758),
            .I(N__22753));
    Span4Mux_h I__4195 (
            .O(N__22753),
            .I(N__22750));
    Span4Mux_h I__4194 (
            .O(N__22750),
            .I(N__22747));
    Odrv4 I__4193 (
            .O(N__22747),
            .I(\this_spr_ram.mem_WE_10 ));
    InMux I__4192 (
            .O(N__22744),
            .I(N__22739));
    InMux I__4191 (
            .O(N__22743),
            .I(N__22736));
    InMux I__4190 (
            .O(N__22742),
            .I(N__22730));
    LocalMux I__4189 (
            .O(N__22739),
            .I(N__22726));
    LocalMux I__4188 (
            .O(N__22736),
            .I(N__22723));
    InMux I__4187 (
            .O(N__22735),
            .I(N__22720));
    InMux I__4186 (
            .O(N__22734),
            .I(N__22717));
    InMux I__4185 (
            .O(N__22733),
            .I(N__22714));
    LocalMux I__4184 (
            .O(N__22730),
            .I(N__22711));
    InMux I__4183 (
            .O(N__22729),
            .I(N__22708));
    Sp12to4 I__4182 (
            .O(N__22726),
            .I(N__22704));
    Span4Mux_h I__4181 (
            .O(N__22723),
            .I(N__22701));
    LocalMux I__4180 (
            .O(N__22720),
            .I(N__22698));
    LocalMux I__4179 (
            .O(N__22717),
            .I(N__22695));
    LocalMux I__4178 (
            .O(N__22714),
            .I(N__22692));
    Span12Mux_h I__4177 (
            .O(N__22711),
            .I(N__22689));
    LocalMux I__4176 (
            .O(N__22708),
            .I(N__22686));
    InMux I__4175 (
            .O(N__22707),
            .I(N__22683));
    Span12Mux_v I__4174 (
            .O(N__22704),
            .I(N__22680));
    Span4Mux_h I__4173 (
            .O(N__22701),
            .I(N__22677));
    Span12Mux_h I__4172 (
            .O(N__22698),
            .I(N__22670));
    Span12Mux_h I__4171 (
            .O(N__22695),
            .I(N__22670));
    Span12Mux_h I__4170 (
            .O(N__22692),
            .I(N__22670));
    Span12Mux_v I__4169 (
            .O(N__22689),
            .I(N__22663));
    Span12Mux_h I__4168 (
            .O(N__22686),
            .I(N__22663));
    LocalMux I__4167 (
            .O(N__22683),
            .I(N__22663));
    Odrv12 I__4166 (
            .O(N__22680),
            .I(M_this_spr_ram_write_data_2));
    Odrv4 I__4165 (
            .O(N__22677),
            .I(M_this_spr_ram_write_data_2));
    Odrv12 I__4164 (
            .O(N__22670),
            .I(M_this_spr_ram_write_data_2));
    Odrv12 I__4163 (
            .O(N__22663),
            .I(M_this_spr_ram_write_data_2));
    CascadeMux I__4162 (
            .O(N__22654),
            .I(N__22651));
    InMux I__4161 (
            .O(N__22651),
            .I(N__22648));
    LocalMux I__4160 (
            .O(N__22648),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ));
    CascadeMux I__4159 (
            .O(N__22645),
            .I(N__22641));
    CascadeMux I__4158 (
            .O(N__22644),
            .I(N__22637));
    InMux I__4157 (
            .O(N__22641),
            .I(N__22634));
    InMux I__4156 (
            .O(N__22640),
            .I(N__22629));
    InMux I__4155 (
            .O(N__22637),
            .I(N__22629));
    LocalMux I__4154 (
            .O(N__22634),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    LocalMux I__4153 (
            .O(N__22629),
            .I(\this_ppu.M_count_qZ0Z_6 ));
    InMux I__4152 (
            .O(N__22624),
            .I(N__22621));
    LocalMux I__4151 (
            .O(N__22621),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ));
    CascadeMux I__4150 (
            .O(N__22618),
            .I(N__22614));
    InMux I__4149 (
            .O(N__22617),
            .I(N__22610));
    InMux I__4148 (
            .O(N__22614),
            .I(N__22605));
    InMux I__4147 (
            .O(N__22613),
            .I(N__22605));
    LocalMux I__4146 (
            .O(N__22610),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    LocalMux I__4145 (
            .O(N__22605),
            .I(\this_ppu.M_count_qZ0Z_3 ));
    IoInMux I__4144 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__4143 (
            .O(N__22597),
            .I(N__22594));
    Odrv4 I__4142 (
            .O(N__22594),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    InMux I__4141 (
            .O(N__22591),
            .I(N__22588));
    LocalMux I__4140 (
            .O(N__22588),
            .I(N__22585));
    Span12Mux_h I__4139 (
            .O(N__22585),
            .I(N__22582));
    Odrv12 I__4138 (
            .O(N__22582),
            .I(\this_spr_ram.mem_out_bus4_3 ));
    InMux I__4137 (
            .O(N__22579),
            .I(N__22576));
    LocalMux I__4136 (
            .O(N__22576),
            .I(N__22573));
    Span12Mux_h I__4135 (
            .O(N__22573),
            .I(N__22570));
    Odrv12 I__4134 (
            .O(N__22570),
            .I(\this_spr_ram.mem_out_bus0_3 ));
    CascadeMux I__4133 (
            .O(N__22567),
            .I(N__22564));
    InMux I__4132 (
            .O(N__22564),
            .I(N__22561));
    LocalMux I__4131 (
            .O(N__22561),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ));
    InMux I__4130 (
            .O(N__22558),
            .I(N__22555));
    LocalMux I__4129 (
            .O(N__22555),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    InMux I__4128 (
            .O(N__22552),
            .I(N__22549));
    LocalMux I__4127 (
            .O(N__22549),
            .I(N__22546));
    Span12Mux_v I__4126 (
            .O(N__22546),
            .I(N__22543));
    Odrv12 I__4125 (
            .O(N__22543),
            .I(\this_spr_ram.mem_out_bus7_3 ));
    InMux I__4124 (
            .O(N__22540),
            .I(N__22537));
    LocalMux I__4123 (
            .O(N__22537),
            .I(N__22534));
    Span4Mux_h I__4122 (
            .O(N__22534),
            .I(N__22531));
    Span4Mux_h I__4121 (
            .O(N__22531),
            .I(N__22528));
    Odrv4 I__4120 (
            .O(N__22528),
            .I(\this_spr_ram.mem_out_bus3_3 ));
    InMux I__4119 (
            .O(N__22525),
            .I(N__22522));
    LocalMux I__4118 (
            .O(N__22522),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ));
    InMux I__4117 (
            .O(N__22519),
            .I(\this_ppu.un1_M_count_q_1_cry_2_s1 ));
    InMux I__4116 (
            .O(N__22516),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1 ));
    InMux I__4115 (
            .O(N__22513),
            .I(\this_ppu.un1_M_count_q_1_cry_4_s1 ));
    InMux I__4114 (
            .O(N__22510),
            .I(\this_ppu.un1_M_count_q_1_cry_5_s1 ));
    InMux I__4113 (
            .O(N__22507),
            .I(\this_ppu.un1_M_count_q_1_cry_6_s1 ));
    InMux I__4112 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__4111 (
            .O(N__22501),
            .I(\this_ppu.M_count_q_RNO_0Z0Z_7 ));
    CascadeMux I__4110 (
            .O(N__22498),
            .I(N__22495));
    InMux I__4109 (
            .O(N__22495),
            .I(N__22492));
    LocalMux I__4108 (
            .O(N__22492),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ));
    CascadeMux I__4107 (
            .O(N__22489),
            .I(N__22485));
    InMux I__4106 (
            .O(N__22488),
            .I(N__22481));
    InMux I__4105 (
            .O(N__22485),
            .I(N__22478));
    InMux I__4104 (
            .O(N__22484),
            .I(N__22475));
    LocalMux I__4103 (
            .O(N__22481),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__4102 (
            .O(N__22478),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    LocalMux I__4101 (
            .O(N__22475),
            .I(\this_ppu.M_count_qZ0Z_2 ));
    CascadeMux I__4100 (
            .O(N__22468),
            .I(\this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_ ));
    CascadeMux I__4099 (
            .O(N__22465),
            .I(N__22462));
    InMux I__4098 (
            .O(N__22462),
            .I(N__22459));
    LocalMux I__4097 (
            .O(N__22459),
            .I(N__22456));
    Odrv4 I__4096 (
            .O(N__22456),
            .I(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ));
    InMux I__4095 (
            .O(N__22453),
            .I(N__22449));
    CascadeMux I__4094 (
            .O(N__22452),
            .I(N__22446));
    LocalMux I__4093 (
            .O(N__22449),
            .I(N__22442));
    InMux I__4092 (
            .O(N__22446),
            .I(N__22439));
    InMux I__4091 (
            .O(N__22445),
            .I(N__22436));
    Odrv4 I__4090 (
            .O(N__22442),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__4089 (
            .O(N__22439),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    LocalMux I__4088 (
            .O(N__22436),
            .I(\this_ppu.M_count_qZ0Z_4 ));
    CascadeMux I__4087 (
            .O(N__22429),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_ ));
    InMux I__4086 (
            .O(N__22426),
            .I(N__22423));
    LocalMux I__4085 (
            .O(N__22423),
            .I(\this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11 ));
    InMux I__4084 (
            .O(N__22420),
            .I(\this_ppu.un1_M_count_q_1_cry_0_s1 ));
    InMux I__4083 (
            .O(N__22417),
            .I(\this_ppu.un1_M_count_q_1_cry_1_s1 ));
    SRMux I__4082 (
            .O(N__22414),
            .I(N__22410));
    SRMux I__4081 (
            .O(N__22413),
            .I(N__22406));
    LocalMux I__4080 (
            .O(N__22410),
            .I(N__22402));
    SRMux I__4079 (
            .O(N__22409),
            .I(N__22399));
    LocalMux I__4078 (
            .O(N__22406),
            .I(N__22396));
    SRMux I__4077 (
            .O(N__22405),
            .I(N__22393));
    Span4Mux_v I__4076 (
            .O(N__22402),
            .I(N__22388));
    LocalMux I__4075 (
            .O(N__22399),
            .I(N__22388));
    Span4Mux_v I__4074 (
            .O(N__22396),
            .I(N__22385));
    LocalMux I__4073 (
            .O(N__22393),
            .I(N__22382));
    Span4Mux_h I__4072 (
            .O(N__22388),
            .I(N__22379));
    Odrv4 I__4071 (
            .O(N__22385),
            .I(\this_ppu.M_last_q_RNIGL6V4 ));
    Odrv12 I__4070 (
            .O(N__22382),
            .I(\this_ppu.M_last_q_RNIGL6V4 ));
    Odrv4 I__4069 (
            .O(N__22379),
            .I(\this_ppu.M_last_q_RNIGL6V4 ));
    CEMux I__4068 (
            .O(N__22372),
            .I(N__22369));
    LocalMux I__4067 (
            .O(N__22369),
            .I(N__22365));
    CEMux I__4066 (
            .O(N__22368),
            .I(N__22362));
    Span4Mux_v I__4065 (
            .O(N__22365),
            .I(N__22357));
    LocalMux I__4064 (
            .O(N__22362),
            .I(N__22357));
    Span4Mux_h I__4063 (
            .O(N__22357),
            .I(N__22354));
    Span4Mux_h I__4062 (
            .O(N__22354),
            .I(N__22351));
    Odrv4 I__4061 (
            .O(N__22351),
            .I(\this_spr_ram.mem_WE_8 ));
    InMux I__4060 (
            .O(N__22348),
            .I(N__22345));
    LocalMux I__4059 (
            .O(N__22345),
            .I(N__22342));
    Span4Mux_h I__4058 (
            .O(N__22342),
            .I(N__22339));
    Span4Mux_v I__4057 (
            .O(N__22339),
            .I(N__22336));
    Span4Mux_v I__4056 (
            .O(N__22336),
            .I(N__22333));
    Span4Mux_h I__4055 (
            .O(N__22333),
            .I(N__22330));
    Odrv4 I__4054 (
            .O(N__22330),
            .I(M_this_map_ram_read_data_6));
    CascadeMux I__4053 (
            .O(N__22327),
            .I(N__22324));
    InMux I__4052 (
            .O(N__22324),
            .I(N__22320));
    InMux I__4051 (
            .O(N__22323),
            .I(N__22315));
    LocalMux I__4050 (
            .O(N__22320),
            .I(N__22312));
    InMux I__4049 (
            .O(N__22319),
            .I(N__22307));
    InMux I__4048 (
            .O(N__22318),
            .I(N__22307));
    LocalMux I__4047 (
            .O(N__22315),
            .I(N__22304));
    Span4Mux_h I__4046 (
            .O(N__22312),
            .I(N__22299));
    LocalMux I__4045 (
            .O(N__22307),
            .I(N__22299));
    Span4Mux_h I__4044 (
            .O(N__22304),
            .I(N__22296));
    Odrv4 I__4043 (
            .O(N__22299),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    Odrv4 I__4042 (
            .O(N__22296),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    InMux I__4041 (
            .O(N__22291),
            .I(N__22288));
    LocalMux I__4040 (
            .O(N__22288),
            .I(N__22285));
    Odrv4 I__4039 (
            .O(N__22285),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    InMux I__4038 (
            .O(N__22282),
            .I(N__22279));
    LocalMux I__4037 (
            .O(N__22279),
            .I(N__22276));
    Span4Mux_v I__4036 (
            .O(N__22276),
            .I(N__22273));
    Sp12to4 I__4035 (
            .O(N__22273),
            .I(N__22270));
    Span12Mux_h I__4034 (
            .O(N__22270),
            .I(N__22267));
    Odrv12 I__4033 (
            .O(N__22267),
            .I(M_this_map_ram_read_data_5));
    InMux I__4032 (
            .O(N__22264),
            .I(N__22258));
    InMux I__4031 (
            .O(N__22263),
            .I(N__22255));
    InMux I__4030 (
            .O(N__22262),
            .I(N__22251));
    CascadeMux I__4029 (
            .O(N__22261),
            .I(N__22248));
    LocalMux I__4028 (
            .O(N__22258),
            .I(N__22244));
    LocalMux I__4027 (
            .O(N__22255),
            .I(N__22241));
    InMux I__4026 (
            .O(N__22254),
            .I(N__22238));
    LocalMux I__4025 (
            .O(N__22251),
            .I(N__22235));
    InMux I__4024 (
            .O(N__22248),
            .I(N__22230));
    InMux I__4023 (
            .O(N__22247),
            .I(N__22227));
    Span4Mux_v I__4022 (
            .O(N__22244),
            .I(N__22224));
    Span4Mux_h I__4021 (
            .O(N__22241),
            .I(N__22221));
    LocalMux I__4020 (
            .O(N__22238),
            .I(N__22216));
    Span4Mux_h I__4019 (
            .O(N__22235),
            .I(N__22216));
    InMux I__4018 (
            .O(N__22234),
            .I(N__22211));
    InMux I__4017 (
            .O(N__22233),
            .I(N__22211));
    LocalMux I__4016 (
            .O(N__22230),
            .I(N__22208));
    LocalMux I__4015 (
            .O(N__22227),
            .I(N__22205));
    Span4Mux_v I__4014 (
            .O(N__22224),
            .I(N__22202));
    Span4Mux_v I__4013 (
            .O(N__22221),
            .I(N__22199));
    Span4Mux_v I__4012 (
            .O(N__22216),
            .I(N__22196));
    LocalMux I__4011 (
            .O(N__22211),
            .I(N__22193));
    Span4Mux_v I__4010 (
            .O(N__22208),
            .I(N__22188));
    Span4Mux_h I__4009 (
            .O(N__22205),
            .I(N__22188));
    Odrv4 I__4008 (
            .O(N__22202),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__4007 (
            .O(N__22199),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__4006 (
            .O(N__22196),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv12 I__4005 (
            .O(N__22193),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__4004 (
            .O(N__22188),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    CEMux I__4003 (
            .O(N__22177),
            .I(N__22174));
    LocalMux I__4002 (
            .O(N__22174),
            .I(N__22170));
    InMux I__4001 (
            .O(N__22173),
            .I(N__22167));
    Span4Mux_v I__4000 (
            .O(N__22170),
            .I(N__22154));
    LocalMux I__3999 (
            .O(N__22167),
            .I(N__22154));
    InMux I__3998 (
            .O(N__22166),
            .I(N__22151));
    InMux I__3997 (
            .O(N__22165),
            .I(N__22146));
    InMux I__3996 (
            .O(N__22164),
            .I(N__22146));
    InMux I__3995 (
            .O(N__22163),
            .I(N__22143));
    InMux I__3994 (
            .O(N__22162),
            .I(N__22140));
    InMux I__3993 (
            .O(N__22161),
            .I(N__22137));
    CascadeMux I__3992 (
            .O(N__22160),
            .I(N__22132));
    CEMux I__3991 (
            .O(N__22159),
            .I(N__22129));
    Span4Mux_h I__3990 (
            .O(N__22154),
            .I(N__22124));
    LocalMux I__3989 (
            .O(N__22151),
            .I(N__22124));
    LocalMux I__3988 (
            .O(N__22146),
            .I(N__22119));
    LocalMux I__3987 (
            .O(N__22143),
            .I(N__22119));
    LocalMux I__3986 (
            .O(N__22140),
            .I(N__22114));
    LocalMux I__3985 (
            .O(N__22137),
            .I(N__22114));
    InMux I__3984 (
            .O(N__22136),
            .I(N__22111));
    InMux I__3983 (
            .O(N__22135),
            .I(N__22108));
    InMux I__3982 (
            .O(N__22132),
            .I(N__22105));
    LocalMux I__3981 (
            .O(N__22129),
            .I(N__22102));
    Span4Mux_h I__3980 (
            .O(N__22124),
            .I(N__22099));
    Span4Mux_v I__3979 (
            .O(N__22119),
            .I(N__22094));
    Span4Mux_h I__3978 (
            .O(N__22114),
            .I(N__22094));
    LocalMux I__3977 (
            .O(N__22111),
            .I(N__22087));
    LocalMux I__3976 (
            .O(N__22108),
            .I(N__22087));
    LocalMux I__3975 (
            .O(N__22105),
            .I(N__22087));
    Span12Mux_v I__3974 (
            .O(N__22102),
            .I(N__22084));
    Span4Mux_v I__3973 (
            .O(N__22099),
            .I(N__22081));
    Span4Mux_h I__3972 (
            .O(N__22094),
            .I(N__22078));
    Span12Mux_h I__3971 (
            .O(N__22087),
            .I(N__22075));
    Odrv12 I__3970 (
            .O(N__22084),
            .I(M_this_state_d_0_sqmuxa));
    Odrv4 I__3969 (
            .O(N__22081),
            .I(M_this_state_d_0_sqmuxa));
    Odrv4 I__3968 (
            .O(N__22078),
            .I(M_this_state_d_0_sqmuxa));
    Odrv12 I__3967 (
            .O(N__22075),
            .I(M_this_state_d_0_sqmuxa));
    InMux I__3966 (
            .O(N__22066),
            .I(N__22063));
    LocalMux I__3965 (
            .O(N__22063),
            .I(N__22060));
    Span4Mux_v I__3964 (
            .O(N__22060),
            .I(N__22057));
    Sp12to4 I__3963 (
            .O(N__22057),
            .I(N__22054));
    Odrv12 I__3962 (
            .O(N__22054),
            .I(\this_spr_ram.mem_out_bus6_1 ));
    InMux I__3961 (
            .O(N__22051),
            .I(N__22048));
    LocalMux I__3960 (
            .O(N__22048),
            .I(N__22045));
    Span4Mux_h I__3959 (
            .O(N__22045),
            .I(N__22042));
    Span4Mux_v I__3958 (
            .O(N__22042),
            .I(N__22039));
    Span4Mux_h I__3957 (
            .O(N__22039),
            .I(N__22036));
    Odrv4 I__3956 (
            .O(N__22036),
            .I(\this_spr_ram.mem_out_bus2_1 ));
    CascadeMux I__3955 (
            .O(N__22033),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_ ));
    InMux I__3954 (
            .O(N__22030),
            .I(N__22027));
    LocalMux I__3953 (
            .O(N__22027),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1 ));
    CEMux I__3952 (
            .O(N__22024),
            .I(N__22021));
    LocalMux I__3951 (
            .O(N__22021),
            .I(N__22017));
    CEMux I__3950 (
            .O(N__22020),
            .I(N__22014));
    Span4Mux_v I__3949 (
            .O(N__22017),
            .I(N__22009));
    LocalMux I__3948 (
            .O(N__22014),
            .I(N__22009));
    Span4Mux_h I__3947 (
            .O(N__22009),
            .I(N__22006));
    Span4Mux_h I__3946 (
            .O(N__22006),
            .I(N__22003));
    Odrv4 I__3945 (
            .O(N__22003),
            .I(\this_spr_ram.mem_WE_6 ));
    InMux I__3944 (
            .O(N__22000),
            .I(N__21997));
    LocalMux I__3943 (
            .O(N__21997),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ));
    CascadeMux I__3942 (
            .O(N__21994),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ));
    InMux I__3941 (
            .O(N__21991),
            .I(N__21987));
    InMux I__3940 (
            .O(N__21990),
            .I(N__21984));
    LocalMux I__3939 (
            .O(N__21987),
            .I(N__21981));
    LocalMux I__3938 (
            .O(N__21984),
            .I(N__21978));
    Odrv4 I__3937 (
            .O(N__21981),
            .I(M_this_spr_ram_read_data_3));
    Odrv4 I__3936 (
            .O(N__21978),
            .I(M_this_spr_ram_read_data_3));
    InMux I__3935 (
            .O(N__21973),
            .I(N__21970));
    LocalMux I__3934 (
            .O(N__21970),
            .I(N__21967));
    Span4Mux_h I__3933 (
            .O(N__21967),
            .I(N__21964));
    Span4Mux_h I__3932 (
            .O(N__21964),
            .I(N__21961));
    Odrv4 I__3931 (
            .O(N__21961),
            .I(\this_spr_ram.mem_out_bus4_1 ));
    InMux I__3930 (
            .O(N__21958),
            .I(N__21955));
    LocalMux I__3929 (
            .O(N__21955),
            .I(N__21952));
    Sp12to4 I__3928 (
            .O(N__21952),
            .I(N__21949));
    Span12Mux_v I__3927 (
            .O(N__21949),
            .I(N__21946));
    Odrv12 I__3926 (
            .O(N__21946),
            .I(\this_spr_ram.mem_out_bus0_1 ));
    InMux I__3925 (
            .O(N__21943),
            .I(N__21940));
    LocalMux I__3924 (
            .O(N__21940),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ));
    InMux I__3923 (
            .O(N__21937),
            .I(N__21934));
    LocalMux I__3922 (
            .O(N__21934),
            .I(\this_ppu.un1_M_haddress_q_c6 ));
    InMux I__3921 (
            .O(N__21931),
            .I(N__21923));
    InMux I__3920 (
            .O(N__21930),
            .I(N__21923));
    InMux I__3919 (
            .O(N__21929),
            .I(N__21920));
    InMux I__3918 (
            .O(N__21928),
            .I(N__21917));
    LocalMux I__3917 (
            .O(N__21923),
            .I(\this_ppu.N_754_0 ));
    LocalMux I__3916 (
            .O(N__21920),
            .I(\this_ppu.N_754_0 ));
    LocalMux I__3915 (
            .O(N__21917),
            .I(\this_ppu.N_754_0 ));
    InMux I__3914 (
            .O(N__21910),
            .I(N__21906));
    InMux I__3913 (
            .O(N__21909),
            .I(N__21903));
    LocalMux I__3912 (
            .O(N__21906),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    LocalMux I__3911 (
            .O(N__21903),
            .I(\this_ppu.un1_M_haddress_q_c2 ));
    InMux I__3910 (
            .O(N__21898),
            .I(N__21895));
    LocalMux I__3909 (
            .O(N__21895),
            .I(\this_ppu.M_state_qZ0Z_8 ));
    InMux I__3908 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__3907 (
            .O(N__21889),
            .I(N__21886));
    Span4Mux_v I__3906 (
            .O(N__21886),
            .I(N__21883));
    Sp12to4 I__3905 (
            .O(N__21883),
            .I(N__21880));
    Odrv12 I__3904 (
            .O(N__21880),
            .I(\this_spr_ram.mem_out_bus6_3 ));
    InMux I__3903 (
            .O(N__21877),
            .I(N__21874));
    LocalMux I__3902 (
            .O(N__21874),
            .I(N__21871));
    Span4Mux_v I__3901 (
            .O(N__21871),
            .I(N__21868));
    Span4Mux_h I__3900 (
            .O(N__21868),
            .I(N__21865));
    Span4Mux_h I__3899 (
            .O(N__21865),
            .I(N__21862));
    Odrv4 I__3898 (
            .O(N__21862),
            .I(\this_spr_ram.mem_out_bus2_3 ));
    InMux I__3897 (
            .O(N__21859),
            .I(N__21856));
    LocalMux I__3896 (
            .O(N__21856),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ));
    InMux I__3895 (
            .O(N__21853),
            .I(N__21850));
    LocalMux I__3894 (
            .O(N__21850),
            .I(N__21846));
    InMux I__3893 (
            .O(N__21849),
            .I(N__21843));
    Odrv4 I__3892 (
            .O(N__21846),
            .I(M_this_spr_ram_read_data_1));
    LocalMux I__3891 (
            .O(N__21843),
            .I(M_this_spr_ram_read_data_1));
    CascadeMux I__3890 (
            .O(N__21838),
            .I(\this_ppu.un1_M_haddress_q_c3_cascade_ ));
    CascadeMux I__3889 (
            .O(N__21835),
            .I(\this_ppu.un1_M_haddress_q_c6_cascade_ ));
    InMux I__3888 (
            .O(N__21832),
            .I(N__21829));
    LocalMux I__3887 (
            .O(N__21829),
            .I(\this_ppu.un1_M_haddress_q_c3 ));
    InMux I__3886 (
            .O(N__21826),
            .I(N__21823));
    LocalMux I__3885 (
            .O(N__21823),
            .I(N__21820));
    Span4Mux_v I__3884 (
            .O(N__21820),
            .I(N__21817));
    Sp12to4 I__3883 (
            .O(N__21817),
            .I(N__21814));
    Span12Mux_h I__3882 (
            .O(N__21814),
            .I(N__21811));
    Odrv12 I__3881 (
            .O(N__21811),
            .I(\this_spr_ram.mem_out_bus7_1 ));
    InMux I__3880 (
            .O(N__21808),
            .I(N__21805));
    LocalMux I__3879 (
            .O(N__21805),
            .I(N__21802));
    Span4Mux_h I__3878 (
            .O(N__21802),
            .I(N__21799));
    Span4Mux_h I__3877 (
            .O(N__21799),
            .I(N__21796));
    Odrv4 I__3876 (
            .O(N__21796),
            .I(\this_spr_ram.mem_out_bus3_1 ));
    InMux I__3875 (
            .O(N__21793),
            .I(N__21790));
    LocalMux I__3874 (
            .O(N__21790),
            .I(N__21787));
    Span4Mux_h I__3873 (
            .O(N__21787),
            .I(N__21784));
    Span4Mux_h I__3872 (
            .O(N__21784),
            .I(N__21781));
    Span4Mux_h I__3871 (
            .O(N__21781),
            .I(N__21778));
    Odrv4 I__3870 (
            .O(N__21778),
            .I(\this_spr_ram.mem_out_bus6_0 ));
    InMux I__3869 (
            .O(N__21775),
            .I(N__21772));
    LocalMux I__3868 (
            .O(N__21772),
            .I(N__21769));
    Span4Mux_h I__3867 (
            .O(N__21769),
            .I(N__21766));
    Span4Mux_v I__3866 (
            .O(N__21766),
            .I(N__21763));
    Span4Mux_h I__3865 (
            .O(N__21763),
            .I(N__21760));
    Odrv4 I__3864 (
            .O(N__21760),
            .I(\this_spr_ram.mem_out_bus2_0 ));
    CascadeMux I__3863 (
            .O(N__21757),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ));
    InMux I__3862 (
            .O(N__21754),
            .I(N__21751));
    LocalMux I__3861 (
            .O(N__21751),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ));
    InMux I__3860 (
            .O(N__21748),
            .I(N__21745));
    LocalMux I__3859 (
            .O(N__21745),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__3858 (
            .O(N__21742),
            .I(N__21739));
    LocalMux I__3857 (
            .O(N__21739),
            .I(N__21736));
    Span12Mux_h I__3856 (
            .O(N__21736),
            .I(N__21733));
    Odrv12 I__3855 (
            .O(N__21733),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__3854 (
            .O(N__21730),
            .I(N__21727));
    LocalMux I__3853 (
            .O(N__21727),
            .I(N__21724));
    Span12Mux_v I__3852 (
            .O(N__21724),
            .I(N__21721));
    Span12Mux_h I__3851 (
            .O(N__21721),
            .I(N__21718));
    Odrv12 I__3850 (
            .O(N__21718),
            .I(\this_ppu.oam_cache.mem_2 ));
    InMux I__3849 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__3848 (
            .O(N__21712),
            .I(N__21709));
    Odrv12 I__3847 (
            .O(N__21709),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2 ));
    InMux I__3846 (
            .O(N__21706),
            .I(N__21703));
    LocalMux I__3845 (
            .O(N__21703),
            .I(N__21700));
    Odrv12 I__3844 (
            .O(N__21700),
            .I(M_this_map_ram_write_data_6));
    InMux I__3843 (
            .O(N__21697),
            .I(N__21694));
    LocalMux I__3842 (
            .O(N__21694),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ));
    InMux I__3841 (
            .O(N__21691),
            .I(N__21688));
    LocalMux I__3840 (
            .O(N__21688),
            .I(N__21685));
    Span4Mux_h I__3839 (
            .O(N__21685),
            .I(N__21682));
    Span4Mux_h I__3838 (
            .O(N__21682),
            .I(N__21679));
    Span4Mux_h I__3837 (
            .O(N__21679),
            .I(N__21676));
    Span4Mux_v I__3836 (
            .O(N__21676),
            .I(N__21673));
    Odrv4 I__3835 (
            .O(N__21673),
            .I(\this_spr_ram.mem_out_bus7_2 ));
    InMux I__3834 (
            .O(N__21670),
            .I(N__21667));
    LocalMux I__3833 (
            .O(N__21667),
            .I(N__21664));
    Span4Mux_h I__3832 (
            .O(N__21664),
            .I(N__21661));
    Span4Mux_h I__3831 (
            .O(N__21661),
            .I(N__21658));
    Odrv4 I__3830 (
            .O(N__21658),
            .I(\this_spr_ram.mem_out_bus3_2 ));
    CascadeMux I__3829 (
            .O(N__21655),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_ ));
    InMux I__3828 (
            .O(N__21652),
            .I(N__21649));
    LocalMux I__3827 (
            .O(N__21649),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2 ));
    InMux I__3826 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__3825 (
            .O(N__21643),
            .I(N__21640));
    Odrv4 I__3824 (
            .O(N__21640),
            .I(M_this_spr_ram_read_data_2));
    CascadeMux I__3823 (
            .O(N__21637),
            .I(M_this_spr_ram_read_data_2_cascade_));
    InMux I__3822 (
            .O(N__21634),
            .I(N__21631));
    LocalMux I__3821 (
            .O(N__21631),
            .I(N__21628));
    Span4Mux_h I__3820 (
            .O(N__21628),
            .I(N__21625));
    Span4Mux_h I__3819 (
            .O(N__21625),
            .I(N__21622));
    Span4Mux_h I__3818 (
            .O(N__21622),
            .I(N__21619));
    Odrv4 I__3817 (
            .O(N__21619),
            .I(\this_spr_ram.mem_out_bus6_2 ));
    InMux I__3816 (
            .O(N__21616),
            .I(N__21613));
    LocalMux I__3815 (
            .O(N__21613),
            .I(N__21610));
    Span4Mux_h I__3814 (
            .O(N__21610),
            .I(N__21607));
    Span4Mux_v I__3813 (
            .O(N__21607),
            .I(N__21604));
    Span4Mux_h I__3812 (
            .O(N__21604),
            .I(N__21601));
    Odrv4 I__3811 (
            .O(N__21601),
            .I(\this_spr_ram.mem_out_bus2_2 ));
    InMux I__3810 (
            .O(N__21598),
            .I(N__21595));
    LocalMux I__3809 (
            .O(N__21595),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ));
    InMux I__3808 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__3807 (
            .O(N__21589),
            .I(N__21586));
    Span4Mux_h I__3806 (
            .O(N__21586),
            .I(N__21583));
    Sp12to4 I__3805 (
            .O(N__21583),
            .I(N__21580));
    Span12Mux_v I__3804 (
            .O(N__21580),
            .I(N__21577));
    Odrv12 I__3803 (
            .O(N__21577),
            .I(\this_spr_ram.mem_out_bus7_0 ));
    InMux I__3802 (
            .O(N__21574),
            .I(N__21571));
    LocalMux I__3801 (
            .O(N__21571),
            .I(N__21568));
    Span4Mux_h I__3800 (
            .O(N__21568),
            .I(N__21565));
    Span4Mux_h I__3799 (
            .O(N__21565),
            .I(N__21562));
    Odrv4 I__3798 (
            .O(N__21562),
            .I(\this_spr_ram.mem_out_bus3_0 ));
    CascadeMux I__3797 (
            .O(N__21559),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_ ));
    InMux I__3796 (
            .O(N__21556),
            .I(N__21552));
    InMux I__3795 (
            .O(N__21555),
            .I(N__21549));
    LocalMux I__3794 (
            .O(N__21552),
            .I(M_this_spr_ram_read_data_0));
    LocalMux I__3793 (
            .O(N__21549),
            .I(M_this_spr_ram_read_data_0));
    InMux I__3792 (
            .O(N__21544),
            .I(N__21541));
    LocalMux I__3791 (
            .O(N__21541),
            .I(N__21538));
    Span4Mux_v I__3790 (
            .O(N__21538),
            .I(N__21535));
    Span4Mux_h I__3789 (
            .O(N__21535),
            .I(N__21532));
    Odrv4 I__3788 (
            .O(N__21532),
            .I(M_this_ppu_vram_data_3));
    InMux I__3787 (
            .O(N__21529),
            .I(N__21524));
    InMux I__3786 (
            .O(N__21528),
            .I(N__21519));
    InMux I__3785 (
            .O(N__21527),
            .I(N__21519));
    LocalMux I__3784 (
            .O(N__21524),
            .I(\this_ppu.N_806 ));
    LocalMux I__3783 (
            .O(N__21519),
            .I(\this_ppu.N_806 ));
    InMux I__3782 (
            .O(N__21514),
            .I(N__21511));
    LocalMux I__3781 (
            .O(N__21511),
            .I(N__21508));
    Span4Mux_v I__3780 (
            .O(N__21508),
            .I(N__21505));
    Span4Mux_h I__3779 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__3778 (
            .O(N__21502),
            .I(M_this_ppu_vram_data_0));
    InMux I__3777 (
            .O(N__21499),
            .I(N__21496));
    LocalMux I__3776 (
            .O(N__21496),
            .I(N__21493));
    Span4Mux_h I__3775 (
            .O(N__21493),
            .I(N__21490));
    Span4Mux_h I__3774 (
            .O(N__21490),
            .I(N__21487));
    Odrv4 I__3773 (
            .O(N__21487),
            .I(\this_spr_ram.mem_out_bus4_0 ));
    InMux I__3772 (
            .O(N__21484),
            .I(N__21481));
    LocalMux I__3771 (
            .O(N__21481),
            .I(N__21478));
    Span12Mux_v I__3770 (
            .O(N__21478),
            .I(N__21475));
    Span12Mux_h I__3769 (
            .O(N__21475),
            .I(N__21472));
    Odrv12 I__3768 (
            .O(N__21472),
            .I(\this_spr_ram.mem_out_bus0_0 ));
    InMux I__3767 (
            .O(N__21469),
            .I(N__21466));
    LocalMux I__3766 (
            .O(N__21466),
            .I(N__21463));
    Span4Mux_h I__3765 (
            .O(N__21463),
            .I(N__21460));
    Span4Mux_h I__3764 (
            .O(N__21460),
            .I(N__21457));
    Odrv4 I__3763 (
            .O(N__21457),
            .I(M_this_map_ram_read_data_2));
    CascadeMux I__3762 (
            .O(N__21454),
            .I(N__21449));
    CascadeMux I__3761 (
            .O(N__21453),
            .I(N__21444));
    CascadeMux I__3760 (
            .O(N__21452),
            .I(N__21441));
    InMux I__3759 (
            .O(N__21449),
            .I(N__21436));
    CascadeMux I__3758 (
            .O(N__21448),
            .I(N__21433));
    CascadeMux I__3757 (
            .O(N__21447),
            .I(N__21430));
    InMux I__3756 (
            .O(N__21444),
            .I(N__21420));
    InMux I__3755 (
            .O(N__21441),
            .I(N__21417));
    CascadeMux I__3754 (
            .O(N__21440),
            .I(N__21414));
    CascadeMux I__3753 (
            .O(N__21439),
            .I(N__21411));
    LocalMux I__3752 (
            .O(N__21436),
            .I(N__21406));
    InMux I__3751 (
            .O(N__21433),
            .I(N__21403));
    InMux I__3750 (
            .O(N__21430),
            .I(N__21400));
    CascadeMux I__3749 (
            .O(N__21429),
            .I(N__21397));
    CascadeMux I__3748 (
            .O(N__21428),
            .I(N__21394));
    CascadeMux I__3747 (
            .O(N__21427),
            .I(N__21391));
    CascadeMux I__3746 (
            .O(N__21426),
            .I(N__21388));
    CascadeMux I__3745 (
            .O(N__21425),
            .I(N__21385));
    CascadeMux I__3744 (
            .O(N__21424),
            .I(N__21382));
    CascadeMux I__3743 (
            .O(N__21423),
            .I(N__21379));
    LocalMux I__3742 (
            .O(N__21420),
            .I(N__21376));
    LocalMux I__3741 (
            .O(N__21417),
            .I(N__21373));
    InMux I__3740 (
            .O(N__21414),
            .I(N__21370));
    InMux I__3739 (
            .O(N__21411),
            .I(N__21367));
    CascadeMux I__3738 (
            .O(N__21410),
            .I(N__21364));
    CascadeMux I__3737 (
            .O(N__21409),
            .I(N__21361));
    Sp12to4 I__3736 (
            .O(N__21406),
            .I(N__21356));
    LocalMux I__3735 (
            .O(N__21403),
            .I(N__21356));
    LocalMux I__3734 (
            .O(N__21400),
            .I(N__21353));
    InMux I__3733 (
            .O(N__21397),
            .I(N__21350));
    InMux I__3732 (
            .O(N__21394),
            .I(N__21347));
    InMux I__3731 (
            .O(N__21391),
            .I(N__21344));
    InMux I__3730 (
            .O(N__21388),
            .I(N__21341));
    InMux I__3729 (
            .O(N__21385),
            .I(N__21338));
    InMux I__3728 (
            .O(N__21382),
            .I(N__21335));
    InMux I__3727 (
            .O(N__21379),
            .I(N__21332));
    Span4Mux_v I__3726 (
            .O(N__21376),
            .I(N__21325));
    Span4Mux_h I__3725 (
            .O(N__21373),
            .I(N__21325));
    LocalMux I__3724 (
            .O(N__21370),
            .I(N__21325));
    LocalMux I__3723 (
            .O(N__21367),
            .I(N__21322));
    InMux I__3722 (
            .O(N__21364),
            .I(N__21319));
    InMux I__3721 (
            .O(N__21361),
            .I(N__21316));
    Span12Mux_s4_v I__3720 (
            .O(N__21356),
            .I(N__21311));
    Span12Mux_s7_h I__3719 (
            .O(N__21353),
            .I(N__21311));
    LocalMux I__3718 (
            .O(N__21350),
            .I(N__21300));
    LocalMux I__3717 (
            .O(N__21347),
            .I(N__21300));
    LocalMux I__3716 (
            .O(N__21344),
            .I(N__21300));
    LocalMux I__3715 (
            .O(N__21341),
            .I(N__21300));
    LocalMux I__3714 (
            .O(N__21338),
            .I(N__21300));
    LocalMux I__3713 (
            .O(N__21335),
            .I(N__21297));
    LocalMux I__3712 (
            .O(N__21332),
            .I(N__21294));
    Span4Mux_v I__3711 (
            .O(N__21325),
            .I(N__21287));
    Span4Mux_h I__3710 (
            .O(N__21322),
            .I(N__21287));
    LocalMux I__3709 (
            .O(N__21319),
            .I(N__21287));
    LocalMux I__3708 (
            .O(N__21316),
            .I(N__21284));
    Span12Mux_h I__3707 (
            .O(N__21311),
            .I(N__21281));
    Span12Mux_v I__3706 (
            .O(N__21300),
            .I(N__21274));
    Span12Mux_v I__3705 (
            .O(N__21297),
            .I(N__21274));
    Span12Mux_s7_h I__3704 (
            .O(N__21294),
            .I(N__21274));
    Span4Mux_v I__3703 (
            .O(N__21287),
            .I(N__21269));
    Span4Mux_h I__3702 (
            .O(N__21284),
            .I(N__21269));
    Span12Mux_v I__3701 (
            .O(N__21281),
            .I(N__21264));
    Span12Mux_h I__3700 (
            .O(N__21274),
            .I(N__21264));
    Span4Mux_h I__3699 (
            .O(N__21269),
            .I(N__21261));
    Odrv12 I__3698 (
            .O(N__21264),
            .I(M_this_ppu_spr_addr_8));
    Odrv4 I__3697 (
            .O(N__21261),
            .I(M_this_ppu_spr_addr_8));
    InMux I__3696 (
            .O(N__21256),
            .I(N__21253));
    LocalMux I__3695 (
            .O(N__21253),
            .I(N__21250));
    Span12Mux_h I__3694 (
            .O(N__21250),
            .I(N__21247));
    Odrv12 I__3693 (
            .O(N__21247),
            .I(M_this_map_ram_read_data_1));
    CascadeMux I__3692 (
            .O(N__21244),
            .I(N__21240));
    CascadeMux I__3691 (
            .O(N__21243),
            .I(N__21237));
    InMux I__3690 (
            .O(N__21240),
            .I(N__21232));
    InMux I__3689 (
            .O(N__21237),
            .I(N__21229));
    CascadeMux I__3688 (
            .O(N__21236),
            .I(N__21226));
    CascadeMux I__3687 (
            .O(N__21235),
            .I(N__21223));
    LocalMux I__3686 (
            .O(N__21232),
            .I(N__21215));
    LocalMux I__3685 (
            .O(N__21229),
            .I(N__21215));
    InMux I__3684 (
            .O(N__21226),
            .I(N__21212));
    InMux I__3683 (
            .O(N__21223),
            .I(N__21209));
    CascadeMux I__3682 (
            .O(N__21222),
            .I(N__21206));
    CascadeMux I__3681 (
            .O(N__21221),
            .I(N__21203));
    CascadeMux I__3680 (
            .O(N__21220),
            .I(N__21197));
    Span4Mux_s3_v I__3679 (
            .O(N__21215),
            .I(N__21189));
    LocalMux I__3678 (
            .O(N__21212),
            .I(N__21189));
    LocalMux I__3677 (
            .O(N__21209),
            .I(N__21189));
    InMux I__3676 (
            .O(N__21206),
            .I(N__21186));
    InMux I__3675 (
            .O(N__21203),
            .I(N__21183));
    CascadeMux I__3674 (
            .O(N__21202),
            .I(N__21180));
    CascadeMux I__3673 (
            .O(N__21201),
            .I(N__21177));
    CascadeMux I__3672 (
            .O(N__21200),
            .I(N__21172));
    InMux I__3671 (
            .O(N__21197),
            .I(N__21168));
    CascadeMux I__3670 (
            .O(N__21196),
            .I(N__21165));
    Span4Mux_v I__3669 (
            .O(N__21189),
            .I(N__21159));
    LocalMux I__3668 (
            .O(N__21186),
            .I(N__21159));
    LocalMux I__3667 (
            .O(N__21183),
            .I(N__21156));
    InMux I__3666 (
            .O(N__21180),
            .I(N__21153));
    InMux I__3665 (
            .O(N__21177),
            .I(N__21150));
    CascadeMux I__3664 (
            .O(N__21176),
            .I(N__21147));
    CascadeMux I__3663 (
            .O(N__21175),
            .I(N__21144));
    InMux I__3662 (
            .O(N__21172),
            .I(N__21141));
    CascadeMux I__3661 (
            .O(N__21171),
            .I(N__21138));
    LocalMux I__3660 (
            .O(N__21168),
            .I(N__21135));
    InMux I__3659 (
            .O(N__21165),
            .I(N__21132));
    CascadeMux I__3658 (
            .O(N__21164),
            .I(N__21129));
    Span4Mux_v I__3657 (
            .O(N__21159),
            .I(N__21119));
    Span4Mux_v I__3656 (
            .O(N__21156),
            .I(N__21119));
    LocalMux I__3655 (
            .O(N__21153),
            .I(N__21119));
    LocalMux I__3654 (
            .O(N__21150),
            .I(N__21119));
    InMux I__3653 (
            .O(N__21147),
            .I(N__21116));
    InMux I__3652 (
            .O(N__21144),
            .I(N__21113));
    LocalMux I__3651 (
            .O(N__21141),
            .I(N__21110));
    InMux I__3650 (
            .O(N__21138),
            .I(N__21107));
    Span4Mux_h I__3649 (
            .O(N__21135),
            .I(N__21102));
    LocalMux I__3648 (
            .O(N__21132),
            .I(N__21102));
    InMux I__3647 (
            .O(N__21129),
            .I(N__21099));
    CascadeMux I__3646 (
            .O(N__21128),
            .I(N__21096));
    Span4Mux_v I__3645 (
            .O(N__21119),
            .I(N__21089));
    LocalMux I__3644 (
            .O(N__21116),
            .I(N__21089));
    LocalMux I__3643 (
            .O(N__21113),
            .I(N__21089));
    Span4Mux_h I__3642 (
            .O(N__21110),
            .I(N__21084));
    LocalMux I__3641 (
            .O(N__21107),
            .I(N__21084));
    Span4Mux_v I__3640 (
            .O(N__21102),
            .I(N__21079));
    LocalMux I__3639 (
            .O(N__21099),
            .I(N__21079));
    InMux I__3638 (
            .O(N__21096),
            .I(N__21076));
    Span4Mux_v I__3637 (
            .O(N__21089),
            .I(N__21073));
    Span4Mux_v I__3636 (
            .O(N__21084),
            .I(N__21066));
    Span4Mux_v I__3635 (
            .O(N__21079),
            .I(N__21066));
    LocalMux I__3634 (
            .O(N__21076),
            .I(N__21066));
    Span4Mux_h I__3633 (
            .O(N__21073),
            .I(N__21063));
    Span4Mux_v I__3632 (
            .O(N__21066),
            .I(N__21060));
    Span4Mux_h I__3631 (
            .O(N__21063),
            .I(N__21057));
    Span4Mux_h I__3630 (
            .O(N__21060),
            .I(N__21054));
    Odrv4 I__3629 (
            .O(N__21057),
            .I(M_this_ppu_spr_addr_7));
    Odrv4 I__3628 (
            .O(N__21054),
            .I(M_this_ppu_spr_addr_7));
    InMux I__3627 (
            .O(N__21049),
            .I(N__21046));
    LocalMux I__3626 (
            .O(N__21046),
            .I(N__21043));
    Span4Mux_h I__3625 (
            .O(N__21043),
            .I(N__21040));
    Span4Mux_h I__3624 (
            .O(N__21040),
            .I(N__21037));
    Odrv4 I__3623 (
            .O(N__21037),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__3622 (
            .O(N__21034),
            .I(N__21031));
    InMux I__3621 (
            .O(N__21031),
            .I(N__21026));
    CascadeMux I__3620 (
            .O(N__21030),
            .I(N__21023));
    CascadeMux I__3619 (
            .O(N__21029),
            .I(N__21020));
    LocalMux I__3618 (
            .O(N__21026),
            .I(N__21005));
    InMux I__3617 (
            .O(N__21023),
            .I(N__21002));
    InMux I__3616 (
            .O(N__21020),
            .I(N__20999));
    CascadeMux I__3615 (
            .O(N__21019),
            .I(N__20996));
    CascadeMux I__3614 (
            .O(N__21018),
            .I(N__20993));
    CascadeMux I__3613 (
            .O(N__21017),
            .I(N__20989));
    CascadeMux I__3612 (
            .O(N__21016),
            .I(N__20986));
    CascadeMux I__3611 (
            .O(N__21015),
            .I(N__20983));
    CascadeMux I__3610 (
            .O(N__21014),
            .I(N__20980));
    CascadeMux I__3609 (
            .O(N__21013),
            .I(N__20977));
    CascadeMux I__3608 (
            .O(N__21012),
            .I(N__20974));
    CascadeMux I__3607 (
            .O(N__21011),
            .I(N__20971));
    CascadeMux I__3606 (
            .O(N__21010),
            .I(N__20968));
    CascadeMux I__3605 (
            .O(N__21009),
            .I(N__20965));
    CascadeMux I__3604 (
            .O(N__21008),
            .I(N__20962));
    Span4Mux_v I__3603 (
            .O(N__21005),
            .I(N__20955));
    LocalMux I__3602 (
            .O(N__21002),
            .I(N__20955));
    LocalMux I__3601 (
            .O(N__20999),
            .I(N__20955));
    InMux I__3600 (
            .O(N__20996),
            .I(N__20952));
    InMux I__3599 (
            .O(N__20993),
            .I(N__20949));
    CascadeMux I__3598 (
            .O(N__20992),
            .I(N__20946));
    InMux I__3597 (
            .O(N__20989),
            .I(N__20943));
    InMux I__3596 (
            .O(N__20986),
            .I(N__20940));
    InMux I__3595 (
            .O(N__20983),
            .I(N__20937));
    InMux I__3594 (
            .O(N__20980),
            .I(N__20934));
    InMux I__3593 (
            .O(N__20977),
            .I(N__20931));
    InMux I__3592 (
            .O(N__20974),
            .I(N__20928));
    InMux I__3591 (
            .O(N__20971),
            .I(N__20925));
    InMux I__3590 (
            .O(N__20968),
            .I(N__20922));
    InMux I__3589 (
            .O(N__20965),
            .I(N__20919));
    InMux I__3588 (
            .O(N__20962),
            .I(N__20916));
    Span4Mux_v I__3587 (
            .O(N__20955),
            .I(N__20909));
    LocalMux I__3586 (
            .O(N__20952),
            .I(N__20909));
    LocalMux I__3585 (
            .O(N__20949),
            .I(N__20909));
    InMux I__3584 (
            .O(N__20946),
            .I(N__20906));
    LocalMux I__3583 (
            .O(N__20943),
            .I(N__20893));
    LocalMux I__3582 (
            .O(N__20940),
            .I(N__20893));
    LocalMux I__3581 (
            .O(N__20937),
            .I(N__20893));
    LocalMux I__3580 (
            .O(N__20934),
            .I(N__20893));
    LocalMux I__3579 (
            .O(N__20931),
            .I(N__20893));
    LocalMux I__3578 (
            .O(N__20928),
            .I(N__20893));
    LocalMux I__3577 (
            .O(N__20925),
            .I(N__20884));
    LocalMux I__3576 (
            .O(N__20922),
            .I(N__20884));
    LocalMux I__3575 (
            .O(N__20919),
            .I(N__20884));
    LocalMux I__3574 (
            .O(N__20916),
            .I(N__20884));
    Span4Mux_v I__3573 (
            .O(N__20909),
            .I(N__20879));
    LocalMux I__3572 (
            .O(N__20906),
            .I(N__20879));
    Span12Mux_s11_v I__3571 (
            .O(N__20893),
            .I(N__20876));
    Span12Mux_v I__3570 (
            .O(N__20884),
            .I(N__20873));
    Span4Mux_v I__3569 (
            .O(N__20879),
            .I(N__20870));
    Span12Mux_h I__3568 (
            .O(N__20876),
            .I(N__20865));
    Span12Mux_h I__3567 (
            .O(N__20873),
            .I(N__20865));
    Span4Mux_h I__3566 (
            .O(N__20870),
            .I(N__20862));
    Odrv12 I__3565 (
            .O(N__20865),
            .I(M_this_ppu_spr_addr_9));
    Odrv4 I__3564 (
            .O(N__20862),
            .I(M_this_ppu_spr_addr_9));
    InMux I__3563 (
            .O(N__20857),
            .I(N__20854));
    LocalMux I__3562 (
            .O(N__20854),
            .I(N__20851));
    Span4Mux_h I__3561 (
            .O(N__20851),
            .I(N__20848));
    Span4Mux_v I__3560 (
            .O(N__20848),
            .I(N__20845));
    Odrv4 I__3559 (
            .O(N__20845),
            .I(M_this_map_ram_read_data_4));
    CascadeMux I__3558 (
            .O(N__20842),
            .I(N__20828));
    CascadeMux I__3557 (
            .O(N__20841),
            .I(N__20825));
    CascadeMux I__3556 (
            .O(N__20840),
            .I(N__20822));
    CascadeMux I__3555 (
            .O(N__20839),
            .I(N__20819));
    CascadeMux I__3554 (
            .O(N__20838),
            .I(N__20816));
    CascadeMux I__3553 (
            .O(N__20837),
            .I(N__20812));
    CascadeMux I__3552 (
            .O(N__20836),
            .I(N__20809));
    CascadeMux I__3551 (
            .O(N__20835),
            .I(N__20806));
    CascadeMux I__3550 (
            .O(N__20834),
            .I(N__20802));
    CascadeMux I__3549 (
            .O(N__20833),
            .I(N__20799));
    CascadeMux I__3548 (
            .O(N__20832),
            .I(N__20796));
    CascadeMux I__3547 (
            .O(N__20831),
            .I(N__20793));
    InMux I__3546 (
            .O(N__20828),
            .I(N__20790));
    InMux I__3545 (
            .O(N__20825),
            .I(N__20787));
    InMux I__3544 (
            .O(N__20822),
            .I(N__20784));
    InMux I__3543 (
            .O(N__20819),
            .I(N__20781));
    InMux I__3542 (
            .O(N__20816),
            .I(N__20776));
    CascadeMux I__3541 (
            .O(N__20815),
            .I(N__20773));
    InMux I__3540 (
            .O(N__20812),
            .I(N__20770));
    InMux I__3539 (
            .O(N__20809),
            .I(N__20767));
    InMux I__3538 (
            .O(N__20806),
            .I(N__20764));
    CascadeMux I__3537 (
            .O(N__20805),
            .I(N__20761));
    InMux I__3536 (
            .O(N__20802),
            .I(N__20758));
    InMux I__3535 (
            .O(N__20799),
            .I(N__20755));
    InMux I__3534 (
            .O(N__20796),
            .I(N__20752));
    InMux I__3533 (
            .O(N__20793),
            .I(N__20749));
    LocalMux I__3532 (
            .O(N__20790),
            .I(N__20744));
    LocalMux I__3531 (
            .O(N__20787),
            .I(N__20744));
    LocalMux I__3530 (
            .O(N__20784),
            .I(N__20739));
    LocalMux I__3529 (
            .O(N__20781),
            .I(N__20739));
    CascadeMux I__3528 (
            .O(N__20780),
            .I(N__20736));
    CascadeMux I__3527 (
            .O(N__20779),
            .I(N__20733));
    LocalMux I__3526 (
            .O(N__20776),
            .I(N__20730));
    InMux I__3525 (
            .O(N__20773),
            .I(N__20727));
    LocalMux I__3524 (
            .O(N__20770),
            .I(N__20722));
    LocalMux I__3523 (
            .O(N__20767),
            .I(N__20722));
    LocalMux I__3522 (
            .O(N__20764),
            .I(N__20719));
    InMux I__3521 (
            .O(N__20761),
            .I(N__20716));
    LocalMux I__3520 (
            .O(N__20758),
            .I(N__20711));
    LocalMux I__3519 (
            .O(N__20755),
            .I(N__20711));
    LocalMux I__3518 (
            .O(N__20752),
            .I(N__20708));
    LocalMux I__3517 (
            .O(N__20749),
            .I(N__20705));
    Span4Mux_v I__3516 (
            .O(N__20744),
            .I(N__20700));
    Span4Mux_v I__3515 (
            .O(N__20739),
            .I(N__20700));
    InMux I__3514 (
            .O(N__20736),
            .I(N__20697));
    InMux I__3513 (
            .O(N__20733),
            .I(N__20694));
    Span4Mux_v I__3512 (
            .O(N__20730),
            .I(N__20689));
    LocalMux I__3511 (
            .O(N__20727),
            .I(N__20689));
    Span4Mux_v I__3510 (
            .O(N__20722),
            .I(N__20684));
    Span4Mux_v I__3509 (
            .O(N__20719),
            .I(N__20684));
    LocalMux I__3508 (
            .O(N__20716),
            .I(N__20679));
    Span4Mux_v I__3507 (
            .O(N__20711),
            .I(N__20679));
    Span4Mux_s1_v I__3506 (
            .O(N__20708),
            .I(N__20674));
    Span4Mux_v I__3505 (
            .O(N__20705),
            .I(N__20674));
    Sp12to4 I__3504 (
            .O(N__20700),
            .I(N__20671));
    LocalMux I__3503 (
            .O(N__20697),
            .I(N__20664));
    LocalMux I__3502 (
            .O(N__20694),
            .I(N__20664));
    Sp12to4 I__3501 (
            .O(N__20689),
            .I(N__20664));
    Span4Mux_h I__3500 (
            .O(N__20684),
            .I(N__20659));
    Span4Mux_v I__3499 (
            .O(N__20679),
            .I(N__20659));
    Sp12to4 I__3498 (
            .O(N__20674),
            .I(N__20656));
    Span12Mux_h I__3497 (
            .O(N__20671),
            .I(N__20653));
    Span12Mux_v I__3496 (
            .O(N__20664),
            .I(N__20650));
    Span4Mux_h I__3495 (
            .O(N__20659),
            .I(N__20647));
    Span12Mux_h I__3494 (
            .O(N__20656),
            .I(N__20644));
    Span12Mux_v I__3493 (
            .O(N__20653),
            .I(N__20641));
    Span12Mux_h I__3492 (
            .O(N__20650),
            .I(N__20634));
    Sp12to4 I__3491 (
            .O(N__20647),
            .I(N__20634));
    Span12Mux_v I__3490 (
            .O(N__20644),
            .I(N__20634));
    Odrv12 I__3489 (
            .O(N__20641),
            .I(M_this_ppu_spr_addr_10));
    Odrv12 I__3488 (
            .O(N__20634),
            .I(M_this_ppu_spr_addr_10));
    InMux I__3487 (
            .O(N__20629),
            .I(N__20626));
    LocalMux I__3486 (
            .O(N__20626),
            .I(N__20623));
    Span12Mux_v I__3485 (
            .O(N__20623),
            .I(N__20620));
    Span12Mux_h I__3484 (
            .O(N__20620),
            .I(N__20617));
    Odrv12 I__3483 (
            .O(N__20617),
            .I(\this_ppu.oam_cache.mem_3 ));
    InMux I__3482 (
            .O(N__20614),
            .I(N__20611));
    LocalMux I__3481 (
            .O(N__20611),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_3 ));
    CascadeMux I__3480 (
            .O(N__20608),
            .I(N__20603));
    InMux I__3479 (
            .O(N__20607),
            .I(N__20599));
    InMux I__3478 (
            .O(N__20606),
            .I(N__20596));
    InMux I__3477 (
            .O(N__20603),
            .I(N__20593));
    InMux I__3476 (
            .O(N__20602),
            .I(N__20590));
    LocalMux I__3475 (
            .O(N__20599),
            .I(this_vga_signals_M_lcounter_q_0));
    LocalMux I__3474 (
            .O(N__20596),
            .I(this_vga_signals_M_lcounter_q_0));
    LocalMux I__3473 (
            .O(N__20593),
            .I(this_vga_signals_M_lcounter_q_0));
    LocalMux I__3472 (
            .O(N__20590),
            .I(this_vga_signals_M_lcounter_q_0));
    InMux I__3471 (
            .O(N__20581),
            .I(N__20577));
    InMux I__3470 (
            .O(N__20580),
            .I(N__20574));
    LocalMux I__3469 (
            .O(N__20577),
            .I(N__20571));
    LocalMux I__3468 (
            .O(N__20574),
            .I(N__20568));
    Span4Mux_v I__3467 (
            .O(N__20571),
            .I(N__20565));
    Span4Mux_h I__3466 (
            .O(N__20568),
            .I(N__20562));
    Span4Mux_h I__3465 (
            .O(N__20565),
            .I(N__20557));
    Span4Mux_v I__3464 (
            .O(N__20562),
            .I(N__20557));
    Odrv4 I__3463 (
            .O(N__20557),
            .I(\this_ppu.N_759_0 ));
    CascadeMux I__3462 (
            .O(N__20554),
            .I(N__20548));
    CascadeMux I__3461 (
            .O(N__20553),
            .I(N__20545));
    CascadeMux I__3460 (
            .O(N__20552),
            .I(N__20542));
    CascadeMux I__3459 (
            .O(N__20551),
            .I(N__20539));
    InMux I__3458 (
            .O(N__20548),
            .I(N__20536));
    InMux I__3457 (
            .O(N__20545),
            .I(N__20533));
    InMux I__3456 (
            .O(N__20542),
            .I(N__20530));
    InMux I__3455 (
            .O(N__20539),
            .I(N__20527));
    LocalMux I__3454 (
            .O(N__20536),
            .I(this_vga_signals_M_lcounter_q_1));
    LocalMux I__3453 (
            .O(N__20533),
            .I(this_vga_signals_M_lcounter_q_1));
    LocalMux I__3452 (
            .O(N__20530),
            .I(this_vga_signals_M_lcounter_q_1));
    LocalMux I__3451 (
            .O(N__20527),
            .I(this_vga_signals_M_lcounter_q_1));
    InMux I__3450 (
            .O(N__20518),
            .I(N__20515));
    LocalMux I__3449 (
            .O(N__20515),
            .I(N__20507));
    InMux I__3448 (
            .O(N__20514),
            .I(N__20504));
    InMux I__3447 (
            .O(N__20513),
            .I(N__20501));
    InMux I__3446 (
            .O(N__20512),
            .I(N__20498));
    InMux I__3445 (
            .O(N__20511),
            .I(N__20495));
    InMux I__3444 (
            .O(N__20510),
            .I(N__20492));
    Span4Mux_h I__3443 (
            .O(N__20507),
            .I(N__20485));
    LocalMux I__3442 (
            .O(N__20504),
            .I(N__20485));
    LocalMux I__3441 (
            .O(N__20501),
            .I(N__20485));
    LocalMux I__3440 (
            .O(N__20498),
            .I(N__20480));
    LocalMux I__3439 (
            .O(N__20495),
            .I(N__20475));
    LocalMux I__3438 (
            .O(N__20492),
            .I(N__20470));
    Span4Mux_h I__3437 (
            .O(N__20485),
            .I(N__20467));
    InMux I__3436 (
            .O(N__20484),
            .I(N__20464));
    InMux I__3435 (
            .O(N__20483),
            .I(N__20461));
    Span4Mux_h I__3434 (
            .O(N__20480),
            .I(N__20458));
    CascadeMux I__3433 (
            .O(N__20479),
            .I(N__20455));
    InMux I__3432 (
            .O(N__20478),
            .I(N__20452));
    Span4Mux_h I__3431 (
            .O(N__20475),
            .I(N__20449));
    InMux I__3430 (
            .O(N__20474),
            .I(N__20444));
    InMux I__3429 (
            .O(N__20473),
            .I(N__20444));
    Span4Mux_v I__3428 (
            .O(N__20470),
            .I(N__20440));
    Span4Mux_h I__3427 (
            .O(N__20467),
            .I(N__20437));
    LocalMux I__3426 (
            .O(N__20464),
            .I(N__20430));
    LocalMux I__3425 (
            .O(N__20461),
            .I(N__20430));
    Span4Mux_h I__3424 (
            .O(N__20458),
            .I(N__20430));
    InMux I__3423 (
            .O(N__20455),
            .I(N__20427));
    LocalMux I__3422 (
            .O(N__20452),
            .I(N__20420));
    Span4Mux_h I__3421 (
            .O(N__20449),
            .I(N__20420));
    LocalMux I__3420 (
            .O(N__20444),
            .I(N__20420));
    InMux I__3419 (
            .O(N__20443),
            .I(N__20417));
    Odrv4 I__3418 (
            .O(N__20440),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3417 (
            .O(N__20437),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3416 (
            .O(N__20430),
            .I(this_vga_signals_M_vcounter_q_9));
    LocalMux I__3415 (
            .O(N__20427),
            .I(this_vga_signals_M_vcounter_q_9));
    Odrv4 I__3414 (
            .O(N__20420),
            .I(this_vga_signals_M_vcounter_q_9));
    LocalMux I__3413 (
            .O(N__20417),
            .I(this_vga_signals_M_vcounter_q_9));
    CascadeMux I__3412 (
            .O(N__20404),
            .I(\this_ppu.N_5_4_cascade_ ));
    InMux I__3411 (
            .O(N__20401),
            .I(N__20398));
    LocalMux I__3410 (
            .O(N__20398),
            .I(N__20395));
    Span4Mux_v I__3409 (
            .O(N__20395),
            .I(N__20392));
    Sp12to4 I__3408 (
            .O(N__20392),
            .I(N__20389));
    Span12Mux_h I__3407 (
            .O(N__20389),
            .I(N__20386));
    Odrv12 I__3406 (
            .O(N__20386),
            .I(\this_ppu.oam_cache.mem_0 ));
    InMux I__3405 (
            .O(N__20383),
            .I(N__20380));
    LocalMux I__3404 (
            .O(N__20380),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ));
    InMux I__3403 (
            .O(N__20377),
            .I(N__20374));
    LocalMux I__3402 (
            .O(N__20374),
            .I(N__20371));
    Span4Mux_h I__3401 (
            .O(N__20371),
            .I(N__20368));
    Odrv4 I__3400 (
            .O(N__20368),
            .I(M_this_map_ram_read_data_0));
    CascadeMux I__3399 (
            .O(N__20365),
            .I(N__20359));
    CascadeMux I__3398 (
            .O(N__20364),
            .I(N__20356));
    CascadeMux I__3397 (
            .O(N__20363),
            .I(N__20352));
    CascadeMux I__3396 (
            .O(N__20362),
            .I(N__20347));
    InMux I__3395 (
            .O(N__20359),
            .I(N__20343));
    InMux I__3394 (
            .O(N__20356),
            .I(N__20339));
    CascadeMux I__3393 (
            .O(N__20355),
            .I(N__20336));
    InMux I__3392 (
            .O(N__20352),
            .I(N__20332));
    CascadeMux I__3391 (
            .O(N__20351),
            .I(N__20329));
    CascadeMux I__3390 (
            .O(N__20350),
            .I(N__20326));
    InMux I__3389 (
            .O(N__20347),
            .I(N__20322));
    CascadeMux I__3388 (
            .O(N__20346),
            .I(N__20319));
    LocalMux I__3387 (
            .O(N__20343),
            .I(N__20316));
    CascadeMux I__3386 (
            .O(N__20342),
            .I(N__20313));
    LocalMux I__3385 (
            .O(N__20339),
            .I(N__20309));
    InMux I__3384 (
            .O(N__20336),
            .I(N__20306));
    CascadeMux I__3383 (
            .O(N__20335),
            .I(N__20303));
    LocalMux I__3382 (
            .O(N__20332),
            .I(N__20299));
    InMux I__3381 (
            .O(N__20329),
            .I(N__20296));
    InMux I__3380 (
            .O(N__20326),
            .I(N__20293));
    CascadeMux I__3379 (
            .O(N__20325),
            .I(N__20290));
    LocalMux I__3378 (
            .O(N__20322),
            .I(N__20287));
    InMux I__3377 (
            .O(N__20319),
            .I(N__20284));
    Span4Mux_v I__3376 (
            .O(N__20316),
            .I(N__20281));
    InMux I__3375 (
            .O(N__20313),
            .I(N__20278));
    CascadeMux I__3374 (
            .O(N__20312),
            .I(N__20275));
    Span4Mux_h I__3373 (
            .O(N__20309),
            .I(N__20269));
    LocalMux I__3372 (
            .O(N__20306),
            .I(N__20269));
    InMux I__3371 (
            .O(N__20303),
            .I(N__20266));
    CascadeMux I__3370 (
            .O(N__20302),
            .I(N__20263));
    Span4Mux_h I__3369 (
            .O(N__20299),
            .I(N__20257));
    LocalMux I__3368 (
            .O(N__20296),
            .I(N__20257));
    LocalMux I__3367 (
            .O(N__20293),
            .I(N__20254));
    InMux I__3366 (
            .O(N__20290),
            .I(N__20251));
    Span4Mux_v I__3365 (
            .O(N__20287),
            .I(N__20246));
    LocalMux I__3364 (
            .O(N__20284),
            .I(N__20246));
    Span4Mux_v I__3363 (
            .O(N__20281),
            .I(N__20241));
    LocalMux I__3362 (
            .O(N__20278),
            .I(N__20241));
    InMux I__3361 (
            .O(N__20275),
            .I(N__20238));
    CascadeMux I__3360 (
            .O(N__20274),
            .I(N__20235));
    Span4Mux_v I__3359 (
            .O(N__20269),
            .I(N__20229));
    LocalMux I__3358 (
            .O(N__20266),
            .I(N__20229));
    InMux I__3357 (
            .O(N__20263),
            .I(N__20226));
    CascadeMux I__3356 (
            .O(N__20262),
            .I(N__20223));
    Span4Mux_v I__3355 (
            .O(N__20257),
            .I(N__20218));
    Span4Mux_h I__3354 (
            .O(N__20254),
            .I(N__20218));
    LocalMux I__3353 (
            .O(N__20251),
            .I(N__20215));
    Span4Mux_v I__3352 (
            .O(N__20246),
            .I(N__20208));
    Span4Mux_h I__3351 (
            .O(N__20241),
            .I(N__20208));
    LocalMux I__3350 (
            .O(N__20238),
            .I(N__20208));
    InMux I__3349 (
            .O(N__20235),
            .I(N__20205));
    CascadeMux I__3348 (
            .O(N__20234),
            .I(N__20202));
    Span4Mux_h I__3347 (
            .O(N__20229),
            .I(N__20197));
    LocalMux I__3346 (
            .O(N__20226),
            .I(N__20197));
    InMux I__3345 (
            .O(N__20223),
            .I(N__20194));
    Span4Mux_h I__3344 (
            .O(N__20218),
            .I(N__20191));
    Span12Mux_s8_h I__3343 (
            .O(N__20215),
            .I(N__20188));
    Span4Mux_v I__3342 (
            .O(N__20208),
            .I(N__20185));
    LocalMux I__3341 (
            .O(N__20205),
            .I(N__20182));
    InMux I__3340 (
            .O(N__20202),
            .I(N__20179));
    Span4Mux_v I__3339 (
            .O(N__20197),
            .I(N__20174));
    LocalMux I__3338 (
            .O(N__20194),
            .I(N__20174));
    Span4Mux_h I__3337 (
            .O(N__20191),
            .I(N__20171));
    Span12Mux_h I__3336 (
            .O(N__20188),
            .I(N__20168));
    Sp12to4 I__3335 (
            .O(N__20185),
            .I(N__20163));
    Span12Mux_s8_h I__3334 (
            .O(N__20182),
            .I(N__20163));
    LocalMux I__3333 (
            .O(N__20179),
            .I(N__20160));
    Span4Mux_v I__3332 (
            .O(N__20174),
            .I(N__20157));
    Span4Mux_h I__3331 (
            .O(N__20171),
            .I(N__20154));
    Span12Mux_v I__3330 (
            .O(N__20168),
            .I(N__20147));
    Span12Mux_h I__3329 (
            .O(N__20163),
            .I(N__20147));
    Span12Mux_s11_h I__3328 (
            .O(N__20160),
            .I(N__20147));
    Span4Mux_h I__3327 (
            .O(N__20157),
            .I(N__20144));
    Odrv4 I__3326 (
            .O(N__20154),
            .I(M_this_ppu_spr_addr_6));
    Odrv12 I__3325 (
            .O(N__20147),
            .I(M_this_ppu_spr_addr_6));
    Odrv4 I__3324 (
            .O(N__20144),
            .I(M_this_ppu_spr_addr_6));
    InMux I__3323 (
            .O(N__20137),
            .I(N__20134));
    LocalMux I__3322 (
            .O(N__20134),
            .I(N__20131));
    Span4Mux_v I__3321 (
            .O(N__20131),
            .I(N__20128));
    Span4Mux_h I__3320 (
            .O(N__20128),
            .I(N__20125));
    Odrv4 I__3319 (
            .O(N__20125),
            .I(\this_spr_ram.mem_out_bus4_2 ));
    InMux I__3318 (
            .O(N__20122),
            .I(N__20119));
    LocalMux I__3317 (
            .O(N__20119),
            .I(N__20116));
    Span12Mux_v I__3316 (
            .O(N__20116),
            .I(N__20113));
    Span12Mux_h I__3315 (
            .O(N__20113),
            .I(N__20110));
    Odrv12 I__3314 (
            .O(N__20110),
            .I(\this_spr_ram.mem_out_bus0_2 ));
    CEMux I__3313 (
            .O(N__20107),
            .I(N__20104));
    LocalMux I__3312 (
            .O(N__20104),
            .I(N__20101));
    Span4Mux_h I__3311 (
            .O(N__20101),
            .I(N__20098));
    Span4Mux_h I__3310 (
            .O(N__20098),
            .I(N__20095));
    Odrv4 I__3309 (
            .O(N__20095),
            .I(M_state_q_RNIQER3C_9));
    InMux I__3308 (
            .O(N__20092),
            .I(N__20089));
    LocalMux I__3307 (
            .O(N__20089),
            .I(N__20086));
    Span4Mux_v I__3306 (
            .O(N__20086),
            .I(N__20083));
    Span4Mux_h I__3305 (
            .O(N__20083),
            .I(N__20080));
    Odrv4 I__3304 (
            .O(N__20080),
            .I(M_this_ppu_vram_data_1));
    InMux I__3303 (
            .O(N__20077),
            .I(N__20058));
    InMux I__3302 (
            .O(N__20076),
            .I(N__20058));
    InMux I__3301 (
            .O(N__20075),
            .I(N__20048));
    InMux I__3300 (
            .O(N__20074),
            .I(N__20048));
    InMux I__3299 (
            .O(N__20073),
            .I(N__20048));
    InMux I__3298 (
            .O(N__20072),
            .I(N__20048));
    InMux I__3297 (
            .O(N__20071),
            .I(N__20043));
    InMux I__3296 (
            .O(N__20070),
            .I(N__20043));
    InMux I__3295 (
            .O(N__20069),
            .I(N__20038));
    InMux I__3294 (
            .O(N__20068),
            .I(N__20038));
    InMux I__3293 (
            .O(N__20067),
            .I(N__20031));
    InMux I__3292 (
            .O(N__20066),
            .I(N__20031));
    InMux I__3291 (
            .O(N__20065),
            .I(N__20031));
    InMux I__3290 (
            .O(N__20064),
            .I(N__20026));
    CEMux I__3289 (
            .O(N__20063),
            .I(N__20021));
    LocalMux I__3288 (
            .O(N__20058),
            .I(N__20018));
    InMux I__3287 (
            .O(N__20057),
            .I(N__20015));
    LocalMux I__3286 (
            .O(N__20048),
            .I(N__20012));
    LocalMux I__3285 (
            .O(N__20043),
            .I(N__20007));
    LocalMux I__3284 (
            .O(N__20038),
            .I(N__20007));
    LocalMux I__3283 (
            .O(N__20031),
            .I(N__20003));
    InMux I__3282 (
            .O(N__20030),
            .I(N__20000));
    InMux I__3281 (
            .O(N__20029),
            .I(N__19997));
    LocalMux I__3280 (
            .O(N__20026),
            .I(N__19994));
    InMux I__3279 (
            .O(N__20025),
            .I(N__19991));
    InMux I__3278 (
            .O(N__20024),
            .I(N__19988));
    LocalMux I__3277 (
            .O(N__20021),
            .I(N__19984));
    Span4Mux_h I__3276 (
            .O(N__20018),
            .I(N__19981));
    LocalMux I__3275 (
            .O(N__20015),
            .I(N__19974));
    Span4Mux_v I__3274 (
            .O(N__20012),
            .I(N__19974));
    Span4Mux_h I__3273 (
            .O(N__20007),
            .I(N__19974));
    InMux I__3272 (
            .O(N__20006),
            .I(N__19971));
    Span4Mux_v I__3271 (
            .O(N__20003),
            .I(N__19966));
    LocalMux I__3270 (
            .O(N__20000),
            .I(N__19966));
    LocalMux I__3269 (
            .O(N__19997),
            .I(N__19959));
    Span4Mux_v I__3268 (
            .O(N__19994),
            .I(N__19959));
    LocalMux I__3267 (
            .O(N__19991),
            .I(N__19959));
    LocalMux I__3266 (
            .O(N__19988),
            .I(N__19956));
    InMux I__3265 (
            .O(N__19987),
            .I(N__19952));
    Span4Mux_v I__3264 (
            .O(N__19984),
            .I(N__19947));
    Span4Mux_v I__3263 (
            .O(N__19981),
            .I(N__19947));
    Span4Mux_v I__3262 (
            .O(N__19974),
            .I(N__19944));
    LocalMux I__3261 (
            .O(N__19971),
            .I(N__19941));
    Span4Mux_h I__3260 (
            .O(N__19966),
            .I(N__19938));
    Span4Mux_h I__3259 (
            .O(N__19959),
            .I(N__19935));
    Span4Mux_v I__3258 (
            .O(N__19956),
            .I(N__19932));
    InMux I__3257 (
            .O(N__19955),
            .I(N__19929));
    LocalMux I__3256 (
            .O(N__19952),
            .I(N__19926));
    Span4Mux_v I__3255 (
            .O(N__19947),
            .I(N__19923));
    Span4Mux_h I__3254 (
            .O(N__19944),
            .I(N__19920));
    Span12Mux_v I__3253 (
            .O(N__19941),
            .I(N__19917));
    Span4Mux_v I__3252 (
            .O(N__19938),
            .I(N__19912));
    Span4Mux_h I__3251 (
            .O(N__19935),
            .I(N__19912));
    Span4Mux_v I__3250 (
            .O(N__19932),
            .I(N__19909));
    LocalMux I__3249 (
            .O(N__19929),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv4 I__3248 (
            .O(N__19926),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv4 I__3247 (
            .O(N__19923),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv4 I__3246 (
            .O(N__19920),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv12 I__3245 (
            .O(N__19917),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv4 I__3244 (
            .O(N__19912),
            .I(\this_vga_signals.GZ0Z_406 ));
    Odrv4 I__3243 (
            .O(N__19909),
            .I(\this_vga_signals.GZ0Z_406 ));
    CascadeMux I__3242 (
            .O(N__19894),
            .I(N__19887));
    InMux I__3241 (
            .O(N__19893),
            .I(N__19882));
    InMux I__3240 (
            .O(N__19892),
            .I(N__19882));
    InMux I__3239 (
            .O(N__19891),
            .I(N__19877));
    InMux I__3238 (
            .O(N__19890),
            .I(N__19874));
    InMux I__3237 (
            .O(N__19887),
            .I(N__19871));
    LocalMux I__3236 (
            .O(N__19882),
            .I(N__19867));
    InMux I__3235 (
            .O(N__19881),
            .I(N__19864));
    InMux I__3234 (
            .O(N__19880),
            .I(N__19861));
    LocalMux I__3233 (
            .O(N__19877),
            .I(N__19858));
    LocalMux I__3232 (
            .O(N__19874),
            .I(N__19853));
    LocalMux I__3231 (
            .O(N__19871),
            .I(N__19853));
    InMux I__3230 (
            .O(N__19870),
            .I(N__19850));
    Span4Mux_h I__3229 (
            .O(N__19867),
            .I(N__19843));
    LocalMux I__3228 (
            .O(N__19864),
            .I(N__19843));
    LocalMux I__3227 (
            .O(N__19861),
            .I(N__19840));
    Span4Mux_v I__3226 (
            .O(N__19858),
            .I(N__19836));
    Span4Mux_v I__3225 (
            .O(N__19853),
            .I(N__19833));
    LocalMux I__3224 (
            .O(N__19850),
            .I(N__19830));
    InMux I__3223 (
            .O(N__19849),
            .I(N__19827));
    InMux I__3222 (
            .O(N__19848),
            .I(N__19824));
    Span4Mux_v I__3221 (
            .O(N__19843),
            .I(N__19821));
    Span4Mux_v I__3220 (
            .O(N__19840),
            .I(N__19818));
    InMux I__3219 (
            .O(N__19839),
            .I(N__19815));
    Span4Mux_h I__3218 (
            .O(N__19836),
            .I(N__19808));
    Span4Mux_h I__3217 (
            .O(N__19833),
            .I(N__19808));
    Span4Mux_h I__3216 (
            .O(N__19830),
            .I(N__19808));
    LocalMux I__3215 (
            .O(N__19827),
            .I(\this_vga_signals.N_83_1 ));
    LocalMux I__3214 (
            .O(N__19824),
            .I(\this_vga_signals.N_83_1 ));
    Odrv4 I__3213 (
            .O(N__19821),
            .I(\this_vga_signals.N_83_1 ));
    Odrv4 I__3212 (
            .O(N__19818),
            .I(\this_vga_signals.N_83_1 ));
    LocalMux I__3211 (
            .O(N__19815),
            .I(\this_vga_signals.N_83_1 ));
    Odrv4 I__3210 (
            .O(N__19808),
            .I(\this_vga_signals.N_83_1 ));
    InMux I__3209 (
            .O(N__19795),
            .I(N__19790));
    InMux I__3208 (
            .O(N__19794),
            .I(N__19785));
    InMux I__3207 (
            .O(N__19793),
            .I(N__19785));
    LocalMux I__3206 (
            .O(N__19790),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__3205 (
            .O(N__19785),
            .I(this_pixel_clk_M_counter_q_0));
    InMux I__3204 (
            .O(N__19780),
            .I(N__19777));
    LocalMux I__3203 (
            .O(N__19777),
            .I(N__19774));
    Span4Mux_v I__3202 (
            .O(N__19774),
            .I(N__19771));
    Odrv4 I__3201 (
            .O(N__19771),
            .I(M_this_map_ram_write_data_1));
    InMux I__3200 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__3199 (
            .O(N__19765),
            .I(N__19762));
    Odrv4 I__3198 (
            .O(N__19762),
            .I(M_this_map_ram_write_data_2));
    InMux I__3197 (
            .O(N__19759),
            .I(N__19756));
    LocalMux I__3196 (
            .O(N__19756),
            .I(N__19753));
    Span4Mux_h I__3195 (
            .O(N__19753),
            .I(N__19750));
    Odrv4 I__3194 (
            .O(N__19750),
            .I(M_this_map_ram_write_data_7));
    InMux I__3193 (
            .O(N__19747),
            .I(N__19744));
    LocalMux I__3192 (
            .O(N__19744),
            .I(N__19741));
    Span4Mux_h I__3191 (
            .O(N__19741),
            .I(N__19738));
    Odrv4 I__3190 (
            .O(N__19738),
            .I(M_this_map_ram_write_data_5));
    InMux I__3189 (
            .O(N__19735),
            .I(N__19732));
    LocalMux I__3188 (
            .O(N__19732),
            .I(N__19729));
    Span4Mux_h I__3187 (
            .O(N__19729),
            .I(N__19726));
    Span4Mux_v I__3186 (
            .O(N__19726),
            .I(N__19723));
    Odrv4 I__3185 (
            .O(N__19723),
            .I(M_this_ppu_vram_data_2));
    InMux I__3184 (
            .O(N__19720),
            .I(N__19715));
    InMux I__3183 (
            .O(N__19719),
            .I(N__19712));
    InMux I__3182 (
            .O(N__19718),
            .I(N__19707));
    LocalMux I__3181 (
            .O(N__19715),
            .I(N__19704));
    LocalMux I__3180 (
            .O(N__19712),
            .I(N__19701));
    InMux I__3179 (
            .O(N__19711),
            .I(N__19698));
    CascadeMux I__3178 (
            .O(N__19710),
            .I(N__19695));
    LocalMux I__3177 (
            .O(N__19707),
            .I(N__19692));
    Span4Mux_v I__3176 (
            .O(N__19704),
            .I(N__19689));
    Span4Mux_v I__3175 (
            .O(N__19701),
            .I(N__19684));
    LocalMux I__3174 (
            .O(N__19698),
            .I(N__19684));
    InMux I__3173 (
            .O(N__19695),
            .I(N__19681));
    Span4Mux_v I__3172 (
            .O(N__19692),
            .I(N__19678));
    Span4Mux_h I__3171 (
            .O(N__19689),
            .I(N__19671));
    Span4Mux_v I__3170 (
            .O(N__19684),
            .I(N__19671));
    LocalMux I__3169 (
            .O(N__19681),
            .I(N__19671));
    Odrv4 I__3168 (
            .O(N__19678),
            .I(N_825_0));
    Odrv4 I__3167 (
            .O(N__19671),
            .I(N_825_0));
    InMux I__3166 (
            .O(N__19666),
            .I(N__19660));
    InMux I__3165 (
            .O(N__19665),
            .I(N__19660));
    LocalMux I__3164 (
            .O(N__19660),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__3163 (
            .O(N__19657),
            .I(N__19654));
    LocalMux I__3162 (
            .O(N__19654),
            .I(N__19651));
    Span4Mux_h I__3161 (
            .O(N__19651),
            .I(N__19648));
    Odrv4 I__3160 (
            .O(N__19648),
            .I(M_this_map_ram_write_data_0));
    InMux I__3159 (
            .O(N__19645),
            .I(N__19642));
    LocalMux I__3158 (
            .O(N__19642),
            .I(N__19639));
    Odrv4 I__3157 (
            .O(N__19639),
            .I(M_this_map_ram_write_data_3));
    InMux I__3156 (
            .O(N__19636),
            .I(N__19633));
    LocalMux I__3155 (
            .O(N__19633),
            .I(N__19630));
    Span4Mux_h I__3154 (
            .O(N__19630),
            .I(N__19627));
    Odrv4 I__3153 (
            .O(N__19627),
            .I(M_this_map_ram_write_data_4));
    IoInMux I__3152 (
            .O(N__19624),
            .I(N__19621));
    LocalMux I__3151 (
            .O(N__19621),
            .I(N__19616));
    IoInMux I__3150 (
            .O(N__19620),
            .I(N__19613));
    IoInMux I__3149 (
            .O(N__19619),
            .I(N__19610));
    IoSpan4Mux I__3148 (
            .O(N__19616),
            .I(N__19600));
    LocalMux I__3147 (
            .O(N__19613),
            .I(N__19600));
    LocalMux I__3146 (
            .O(N__19610),
            .I(N__19600));
    IoInMux I__3145 (
            .O(N__19609),
            .I(N__19597));
    IoInMux I__3144 (
            .O(N__19608),
            .I(N__19594));
    IoInMux I__3143 (
            .O(N__19607),
            .I(N__19590));
    IoSpan4Mux I__3142 (
            .O(N__19600),
            .I(N__19580));
    LocalMux I__3141 (
            .O(N__19597),
            .I(N__19580));
    LocalMux I__3140 (
            .O(N__19594),
            .I(N__19577));
    IoInMux I__3139 (
            .O(N__19593),
            .I(N__19574));
    LocalMux I__3138 (
            .O(N__19590),
            .I(N__19571));
    IoInMux I__3137 (
            .O(N__19589),
            .I(N__19568));
    IoInMux I__3136 (
            .O(N__19588),
            .I(N__19565));
    IoInMux I__3135 (
            .O(N__19587),
            .I(N__19561));
    IoInMux I__3134 (
            .O(N__19586),
            .I(N__19558));
    IoInMux I__3133 (
            .O(N__19585),
            .I(N__19555));
    IoSpan4Mux I__3132 (
            .O(N__19580),
            .I(N__19547));
    IoSpan4Mux I__3131 (
            .O(N__19577),
            .I(N__19547));
    LocalMux I__3130 (
            .O(N__19574),
            .I(N__19547));
    IoSpan4Mux I__3129 (
            .O(N__19571),
            .I(N__19540));
    LocalMux I__3128 (
            .O(N__19568),
            .I(N__19540));
    LocalMux I__3127 (
            .O(N__19565),
            .I(N__19540));
    IoInMux I__3126 (
            .O(N__19564),
            .I(N__19537));
    LocalMux I__3125 (
            .O(N__19561),
            .I(N__19531));
    LocalMux I__3124 (
            .O(N__19558),
            .I(N__19531));
    LocalMux I__3123 (
            .O(N__19555),
            .I(N__19528));
    IoInMux I__3122 (
            .O(N__19554),
            .I(N__19525));
    IoSpan4Mux I__3121 (
            .O(N__19547),
            .I(N__19522));
    IoSpan4Mux I__3120 (
            .O(N__19540),
            .I(N__19516));
    LocalMux I__3119 (
            .O(N__19537),
            .I(N__19516));
    IoInMux I__3118 (
            .O(N__19536),
            .I(N__19513));
    IoSpan4Mux I__3117 (
            .O(N__19531),
            .I(N__19510));
    IoSpan4Mux I__3116 (
            .O(N__19528),
            .I(N__19505));
    LocalMux I__3115 (
            .O(N__19525),
            .I(N__19505));
    Span4Mux_s3_v I__3114 (
            .O(N__19522),
            .I(N__19502));
    IoInMux I__3113 (
            .O(N__19521),
            .I(N__19499));
    Sp12to4 I__3112 (
            .O(N__19516),
            .I(N__19494));
    LocalMux I__3111 (
            .O(N__19513),
            .I(N__19494));
    IoSpan4Mux I__3110 (
            .O(N__19510),
            .I(N__19489));
    IoSpan4Mux I__3109 (
            .O(N__19505),
            .I(N__19489));
    Sp12to4 I__3108 (
            .O(N__19502),
            .I(N__19483));
    LocalMux I__3107 (
            .O(N__19499),
            .I(N__19483));
    Span12Mux_s9_h I__3106 (
            .O(N__19494),
            .I(N__19480));
    Sp12to4 I__3105 (
            .O(N__19489),
            .I(N__19477));
    IoInMux I__3104 (
            .O(N__19488),
            .I(N__19474));
    Span12Mux_s10_v I__3103 (
            .O(N__19483),
            .I(N__19471));
    Span12Mux_v I__3102 (
            .O(N__19480),
            .I(N__19466));
    Span12Mux_s9_h I__3101 (
            .O(N__19477),
            .I(N__19466));
    LocalMux I__3100 (
            .O(N__19474),
            .I(N__19463));
    Span12Mux_v I__3099 (
            .O(N__19471),
            .I(N__19460));
    Span12Mux_h I__3098 (
            .O(N__19466),
            .I(N__19455));
    Span12Mux_s10_h I__3097 (
            .O(N__19463),
            .I(N__19455));
    Odrv12 I__3096 (
            .O(N__19460),
            .I(dma_0_i));
    Odrv12 I__3095 (
            .O(N__19455),
            .I(dma_0_i));
    InMux I__3094 (
            .O(N__19450),
            .I(N__19446));
    CascadeMux I__3093 (
            .O(N__19449),
            .I(N__19442));
    LocalMux I__3092 (
            .O(N__19446),
            .I(N__19439));
    InMux I__3091 (
            .O(N__19445),
            .I(N__19436));
    InMux I__3090 (
            .O(N__19442),
            .I(N__19433));
    Span4Mux_h I__3089 (
            .O(N__19439),
            .I(N__19428));
    LocalMux I__3088 (
            .O(N__19436),
            .I(N__19428));
    LocalMux I__3087 (
            .O(N__19433),
            .I(N__19425));
    Span4Mux_v I__3086 (
            .O(N__19428),
            .I(N__19420));
    Span4Mux_v I__3085 (
            .O(N__19425),
            .I(N__19420));
    Odrv4 I__3084 (
            .O(N__19420),
            .I(\this_vga_signals.N_819_0 ));
    CascadeMux I__3083 (
            .O(N__19417),
            .I(\this_vga_signals.N_827_0_cascade_ ));
    InMux I__3082 (
            .O(N__19414),
            .I(N__19411));
    LocalMux I__3081 (
            .O(N__19411),
            .I(\this_vga_signals.N_826_0 ));
    CascadeMux I__3080 (
            .O(N__19408),
            .I(N__19405));
    CascadeBuf I__3079 (
            .O(N__19405),
            .I(N__19402));
    CascadeMux I__3078 (
            .O(N__19402),
            .I(N__19399));
    InMux I__3077 (
            .O(N__19399),
            .I(N__19395));
    InMux I__3076 (
            .O(N__19398),
            .I(N__19392));
    LocalMux I__3075 (
            .O(N__19395),
            .I(N__19389));
    LocalMux I__3074 (
            .O(N__19392),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__3073 (
            .O(N__19389),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__3072 (
            .O(N__19384),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__3071 (
            .O(N__19381),
            .I(N__19378));
    CascadeBuf I__3070 (
            .O(N__19378),
            .I(N__19375));
    CascadeMux I__3069 (
            .O(N__19375),
            .I(N__19372));
    InMux I__3068 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__3067 (
            .O(N__19369),
            .I(N__19365));
    InMux I__3066 (
            .O(N__19368),
            .I(N__19362));
    Span4Mux_h I__3065 (
            .O(N__19365),
            .I(N__19359));
    LocalMux I__3064 (
            .O(N__19362),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__3063 (
            .O(N__19359),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__3062 (
            .O(N__19354),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__3061 (
            .O(N__19351),
            .I(N__19348));
    CascadeBuf I__3060 (
            .O(N__19348),
            .I(N__19345));
    CascadeMux I__3059 (
            .O(N__19345),
            .I(N__19342));
    InMux I__3058 (
            .O(N__19342),
            .I(N__19338));
    InMux I__3057 (
            .O(N__19341),
            .I(N__19335));
    LocalMux I__3056 (
            .O(N__19338),
            .I(N__19332));
    LocalMux I__3055 (
            .O(N__19335),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__3054 (
            .O(N__19332),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__3053 (
            .O(N__19327),
            .I(un1_M_this_map_address_q_cry_4));
    CascadeMux I__3052 (
            .O(N__19324),
            .I(N__19321));
    CascadeBuf I__3051 (
            .O(N__19321),
            .I(N__19318));
    CascadeMux I__3050 (
            .O(N__19318),
            .I(N__19315));
    InMux I__3049 (
            .O(N__19315),
            .I(N__19311));
    InMux I__3048 (
            .O(N__19314),
            .I(N__19308));
    LocalMux I__3047 (
            .O(N__19311),
            .I(N__19305));
    LocalMux I__3046 (
            .O(N__19308),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__3045 (
            .O(N__19305),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__3044 (
            .O(N__19300),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__3043 (
            .O(N__19297),
            .I(N__19294));
    CascadeBuf I__3042 (
            .O(N__19294),
            .I(N__19291));
    CascadeMux I__3041 (
            .O(N__19291),
            .I(N__19288));
    InMux I__3040 (
            .O(N__19288),
            .I(N__19285));
    LocalMux I__3039 (
            .O(N__19285),
            .I(N__19281));
    InMux I__3038 (
            .O(N__19284),
            .I(N__19278));
    Span4Mux_h I__3037 (
            .O(N__19281),
            .I(N__19275));
    LocalMux I__3036 (
            .O(N__19278),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__3035 (
            .O(N__19275),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__3034 (
            .O(N__19270),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__3033 (
            .O(N__19267),
            .I(N__19264));
    CascadeBuf I__3032 (
            .O(N__19264),
            .I(N__19261));
    CascadeMux I__3031 (
            .O(N__19261),
            .I(N__19258));
    InMux I__3030 (
            .O(N__19258),
            .I(N__19255));
    LocalMux I__3029 (
            .O(N__19255),
            .I(N__19251));
    InMux I__3028 (
            .O(N__19254),
            .I(N__19248));
    Span4Mux_h I__3027 (
            .O(N__19251),
            .I(N__19245));
    LocalMux I__3026 (
            .O(N__19248),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__3025 (
            .O(N__19245),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__3024 (
            .O(N__19240),
            .I(bfn_9_22_0_));
    InMux I__3023 (
            .O(N__19237),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__3022 (
            .O(N__19234),
            .I(N__19231));
    CascadeBuf I__3021 (
            .O(N__19231),
            .I(N__19228));
    CascadeMux I__3020 (
            .O(N__19228),
            .I(N__19225));
    InMux I__3019 (
            .O(N__19225),
            .I(N__19221));
    InMux I__3018 (
            .O(N__19224),
            .I(N__19218));
    LocalMux I__3017 (
            .O(N__19221),
            .I(N__19215));
    LocalMux I__3016 (
            .O(N__19218),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__3015 (
            .O(N__19215),
            .I(M_this_map_address_qZ0Z_9));
    IoInMux I__3014 (
            .O(N__19210),
            .I(N__19207));
    LocalMux I__3013 (
            .O(N__19207),
            .I(N__19204));
    IoSpan4Mux I__3012 (
            .O(N__19204),
            .I(N__19201));
    IoSpan4Mux I__3011 (
            .O(N__19201),
            .I(N__19198));
    Span4Mux_s3_v I__3010 (
            .O(N__19198),
            .I(N__19195));
    Odrv4 I__3009 (
            .O(N__19195),
            .I(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ));
    CascadeMux I__3008 (
            .O(N__19192),
            .I(N__19189));
    InMux I__3007 (
            .O(N__19189),
            .I(N__19186));
    LocalMux I__3006 (
            .O(N__19186),
            .I(\this_vga_signals.M_lcounter_q_3_i_o2_0_1 ));
    CascadeMux I__3005 (
            .O(N__19183),
            .I(N__19180));
    InMux I__3004 (
            .O(N__19180),
            .I(N__19175));
    InMux I__3003 (
            .O(N__19179),
            .I(N__19172));
    InMux I__3002 (
            .O(N__19178),
            .I(N__19169));
    LocalMux I__3001 (
            .O(N__19175),
            .I(\this_vga_signals.pixel_clk_i ));
    LocalMux I__3000 (
            .O(N__19172),
            .I(\this_vga_signals.pixel_clk_i ));
    LocalMux I__2999 (
            .O(N__19169),
            .I(\this_vga_signals.pixel_clk_i ));
    CascadeMux I__2998 (
            .O(N__19162),
            .I(\this_vga_signals.N_83_1_cascade_ ));
    InMux I__2997 (
            .O(N__19159),
            .I(N__19153));
    InMux I__2996 (
            .O(N__19158),
            .I(N__19153));
    LocalMux I__2995 (
            .O(N__19153),
            .I(\this_vga_signals.N_2_0 ));
    InMux I__2994 (
            .O(N__19150),
            .I(N__19147));
    LocalMux I__2993 (
            .O(N__19147),
            .I(N__19143));
    InMux I__2992 (
            .O(N__19146),
            .I(N__19140));
    Odrv4 I__2991 (
            .O(N__19143),
            .I(\this_vga_signals.M_pcounter_q_i_2_1 ));
    LocalMux I__2990 (
            .O(N__19140),
            .I(\this_vga_signals.M_pcounter_q_i_2_1 ));
    InMux I__2989 (
            .O(N__19135),
            .I(N__19129));
    InMux I__2988 (
            .O(N__19134),
            .I(N__19126));
    InMux I__2987 (
            .O(N__19133),
            .I(N__19123));
    InMux I__2986 (
            .O(N__19132),
            .I(N__19120));
    LocalMux I__2985 (
            .O(N__19129),
            .I(N__19117));
    LocalMux I__2984 (
            .O(N__19126),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__2983 (
            .O(N__19123),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    LocalMux I__2982 (
            .O(N__19120),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    Odrv4 I__2981 (
            .O(N__19117),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    InMux I__2980 (
            .O(N__19108),
            .I(N__19105));
    LocalMux I__2979 (
            .O(N__19105),
            .I(N__19102));
    Odrv4 I__2978 (
            .O(N__19102),
            .I(\this_vga_signals.M_pcounter_q_0Z0Z_1 ));
    CascadeMux I__2977 (
            .O(N__19099),
            .I(N__19093));
    InMux I__2976 (
            .O(N__19098),
            .I(N__19088));
    InMux I__2975 (
            .O(N__19097),
            .I(N__19085));
    InMux I__2974 (
            .O(N__19096),
            .I(N__19082));
    InMux I__2973 (
            .O(N__19093),
            .I(N__19079));
    InMux I__2972 (
            .O(N__19092),
            .I(N__19076));
    InMux I__2971 (
            .O(N__19091),
            .I(N__19073));
    LocalMux I__2970 (
            .O(N__19088),
            .I(N__19070));
    LocalMux I__2969 (
            .O(N__19085),
            .I(N__19066));
    LocalMux I__2968 (
            .O(N__19082),
            .I(N__19063));
    LocalMux I__2967 (
            .O(N__19079),
            .I(N__19056));
    LocalMux I__2966 (
            .O(N__19076),
            .I(N__19056));
    LocalMux I__2965 (
            .O(N__19073),
            .I(N__19056));
    Span4Mux_v I__2964 (
            .O(N__19070),
            .I(N__19050));
    InMux I__2963 (
            .O(N__19069),
            .I(N__19047));
    Span4Mux_h I__2962 (
            .O(N__19066),
            .I(N__19044));
    Span4Mux_h I__2961 (
            .O(N__19063),
            .I(N__19039));
    Span4Mux_v I__2960 (
            .O(N__19056),
            .I(N__19039));
    InMux I__2959 (
            .O(N__19055),
            .I(N__19036));
    InMux I__2958 (
            .O(N__19054),
            .I(N__19033));
    InMux I__2957 (
            .O(N__19053),
            .I(N__19030));
    Odrv4 I__2956 (
            .O(N__19050),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2955 (
            .O(N__19047),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2954 (
            .O(N__19044),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__2953 (
            .O(N__19039),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2952 (
            .O(N__19036),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2951 (
            .O(N__19033),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__2950 (
            .O(N__19030),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__2949 (
            .O(N__19015),
            .I(N__19010));
    InMux I__2948 (
            .O(N__19014),
            .I(N__19005));
    InMux I__2947 (
            .O(N__19013),
            .I(N__19002));
    LocalMux I__2946 (
            .O(N__19010),
            .I(N__18998));
    InMux I__2945 (
            .O(N__19009),
            .I(N__18992));
    InMux I__2944 (
            .O(N__19008),
            .I(N__18992));
    LocalMux I__2943 (
            .O(N__19005),
            .I(N__18983));
    LocalMux I__2942 (
            .O(N__19002),
            .I(N__18980));
    InMux I__2941 (
            .O(N__19001),
            .I(N__18977));
    Span4Mux_h I__2940 (
            .O(N__18998),
            .I(N__18974));
    InMux I__2939 (
            .O(N__18997),
            .I(N__18971));
    LocalMux I__2938 (
            .O(N__18992),
            .I(N__18968));
    InMux I__2937 (
            .O(N__18991),
            .I(N__18965));
    InMux I__2936 (
            .O(N__18990),
            .I(N__18954));
    InMux I__2935 (
            .O(N__18989),
            .I(N__18954));
    InMux I__2934 (
            .O(N__18988),
            .I(N__18954));
    InMux I__2933 (
            .O(N__18987),
            .I(N__18954));
    InMux I__2932 (
            .O(N__18986),
            .I(N__18954));
    Odrv12 I__2931 (
            .O(N__18983),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2930 (
            .O(N__18980),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2929 (
            .O(N__18977),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2928 (
            .O(N__18974),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2927 (
            .O(N__18971),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__2926 (
            .O(N__18968),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2925 (
            .O(N__18965),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__2924 (
            .O(N__18954),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    InMux I__2923 (
            .O(N__18937),
            .I(N__18933));
    InMux I__2922 (
            .O(N__18936),
            .I(N__18929));
    LocalMux I__2921 (
            .O(N__18933),
            .I(N__18925));
    InMux I__2920 (
            .O(N__18932),
            .I(N__18921));
    LocalMux I__2919 (
            .O(N__18929),
            .I(N__18914));
    InMux I__2918 (
            .O(N__18928),
            .I(N__18911));
    Span4Mux_v I__2917 (
            .O(N__18925),
            .I(N__18908));
    InMux I__2916 (
            .O(N__18924),
            .I(N__18905));
    LocalMux I__2915 (
            .O(N__18921),
            .I(N__18902));
    InMux I__2914 (
            .O(N__18920),
            .I(N__18899));
    InMux I__2913 (
            .O(N__18919),
            .I(N__18896));
    CascadeMux I__2912 (
            .O(N__18918),
            .I(N__18893));
    CascadeMux I__2911 (
            .O(N__18917),
            .I(N__18890));
    Span4Mux_v I__2910 (
            .O(N__18914),
            .I(N__18887));
    LocalMux I__2909 (
            .O(N__18911),
            .I(N__18884));
    Span4Mux_v I__2908 (
            .O(N__18908),
            .I(N__18873));
    LocalMux I__2907 (
            .O(N__18905),
            .I(N__18873));
    Span4Mux_v I__2906 (
            .O(N__18902),
            .I(N__18873));
    LocalMux I__2905 (
            .O(N__18899),
            .I(N__18873));
    LocalMux I__2904 (
            .O(N__18896),
            .I(N__18873));
    InMux I__2903 (
            .O(N__18893),
            .I(N__18870));
    InMux I__2902 (
            .O(N__18890),
            .I(N__18867));
    Odrv4 I__2901 (
            .O(N__18887),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv12 I__2900 (
            .O(N__18884),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__2899 (
            .O(N__18873),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2898 (
            .O(N__18870),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__2897 (
            .O(N__18867),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    CascadeMux I__2896 (
            .O(N__18856),
            .I(\this_vga_signals.N_809_0_cascade_ ));
    CascadeMux I__2895 (
            .O(N__18853),
            .I(N__18850));
    InMux I__2894 (
            .O(N__18850),
            .I(N__18844));
    InMux I__2893 (
            .O(N__18849),
            .I(N__18841));
    InMux I__2892 (
            .O(N__18848),
            .I(N__18836));
    InMux I__2891 (
            .O(N__18847),
            .I(N__18833));
    LocalMux I__2890 (
            .O(N__18844),
            .I(N__18828));
    LocalMux I__2889 (
            .O(N__18841),
            .I(N__18828));
    InMux I__2888 (
            .O(N__18840),
            .I(N__18823));
    InMux I__2887 (
            .O(N__18839),
            .I(N__18823));
    LocalMux I__2886 (
            .O(N__18836),
            .I(N__18820));
    LocalMux I__2885 (
            .O(N__18833),
            .I(N__18816));
    Span4Mux_v I__2884 (
            .O(N__18828),
            .I(N__18810));
    LocalMux I__2883 (
            .O(N__18823),
            .I(N__18810));
    Span4Mux_v I__2882 (
            .O(N__18820),
            .I(N__18806));
    InMux I__2881 (
            .O(N__18819),
            .I(N__18803));
    Span4Mux_h I__2880 (
            .O(N__18816),
            .I(N__18800));
    InMux I__2879 (
            .O(N__18815),
            .I(N__18797));
    Span4Mux_h I__2878 (
            .O(N__18810),
            .I(N__18794));
    InMux I__2877 (
            .O(N__18809),
            .I(N__18791));
    Odrv4 I__2876 (
            .O(N__18806),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2875 (
            .O(N__18803),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2874 (
            .O(N__18800),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2873 (
            .O(N__18797),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__2872 (
            .O(N__18794),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__2871 (
            .O(N__18791),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__2870 (
            .O(N__18778),
            .I(N__18775));
    InMux I__2869 (
            .O(N__18775),
            .I(N__18772));
    LocalMux I__2868 (
            .O(N__18772),
            .I(N__18769));
    Span4Mux_v I__2867 (
            .O(N__18769),
            .I(N__18766));
    Span4Mux_v I__2866 (
            .O(N__18766),
            .I(N__18763));
    Odrv4 I__2865 (
            .O(N__18763),
            .I(N_34_0));
    IoInMux I__2864 (
            .O(N__18760),
            .I(N__18757));
    LocalMux I__2863 (
            .O(N__18757),
            .I(N__18754));
    Span4Mux_s2_h I__2862 (
            .O(N__18754),
            .I(N__18751));
    Span4Mux_v I__2861 (
            .O(N__18751),
            .I(N__18748));
    Span4Mux_h I__2860 (
            .O(N__18748),
            .I(N__18745));
    Odrv4 I__2859 (
            .O(N__18745),
            .I(port_nmib_1_i));
    CascadeMux I__2858 (
            .O(N__18742),
            .I(N__18739));
    CascadeBuf I__2857 (
            .O(N__18739),
            .I(N__18736));
    CascadeMux I__2856 (
            .O(N__18736),
            .I(N__18733));
    InMux I__2855 (
            .O(N__18733),
            .I(N__18730));
    LocalMux I__2854 (
            .O(N__18730),
            .I(N__18726));
    InMux I__2853 (
            .O(N__18729),
            .I(N__18723));
    Span4Mux_v I__2852 (
            .O(N__18726),
            .I(N__18720));
    LocalMux I__2851 (
            .O(N__18723),
            .I(M_this_map_address_qZ0Z_0));
    Odrv4 I__2850 (
            .O(N__18720),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__2849 (
            .O(N__18715),
            .I(N__18712));
    CascadeBuf I__2848 (
            .O(N__18712),
            .I(N__18709));
    CascadeMux I__2847 (
            .O(N__18709),
            .I(N__18706));
    InMux I__2846 (
            .O(N__18706),
            .I(N__18703));
    LocalMux I__2845 (
            .O(N__18703),
            .I(N__18699));
    InMux I__2844 (
            .O(N__18702),
            .I(N__18696));
    Span4Mux_v I__2843 (
            .O(N__18699),
            .I(N__18693));
    LocalMux I__2842 (
            .O(N__18696),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__2841 (
            .O(N__18693),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__2840 (
            .O(N__18688),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__2839 (
            .O(N__18685),
            .I(N__18682));
    CascadeBuf I__2838 (
            .O(N__18682),
            .I(N__18679));
    CascadeMux I__2837 (
            .O(N__18679),
            .I(N__18676));
    InMux I__2836 (
            .O(N__18676),
            .I(N__18673));
    LocalMux I__2835 (
            .O(N__18673),
            .I(N__18669));
    InMux I__2834 (
            .O(N__18672),
            .I(N__18666));
    Span4Mux_h I__2833 (
            .O(N__18669),
            .I(N__18663));
    LocalMux I__2832 (
            .O(N__18666),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__2831 (
            .O(N__18663),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__2830 (
            .O(N__18658),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__2829 (
            .O(N__18655),
            .I(N__18651));
    CascadeMux I__2828 (
            .O(N__18654),
            .I(N__18647));
    InMux I__2827 (
            .O(N__18651),
            .I(N__18641));
    InMux I__2826 (
            .O(N__18650),
            .I(N__18637));
    InMux I__2825 (
            .O(N__18647),
            .I(N__18632));
    InMux I__2824 (
            .O(N__18646),
            .I(N__18632));
    InMux I__2823 (
            .O(N__18645),
            .I(N__18629));
    InMux I__2822 (
            .O(N__18644),
            .I(N__18626));
    LocalMux I__2821 (
            .O(N__18641),
            .I(N__18619));
    InMux I__2820 (
            .O(N__18640),
            .I(N__18616));
    LocalMux I__2819 (
            .O(N__18637),
            .I(N__18613));
    LocalMux I__2818 (
            .O(N__18632),
            .I(N__18608));
    LocalMux I__2817 (
            .O(N__18629),
            .I(N__18608));
    LocalMux I__2816 (
            .O(N__18626),
            .I(N__18604));
    InMux I__2815 (
            .O(N__18625),
            .I(N__18599));
    InMux I__2814 (
            .O(N__18624),
            .I(N__18599));
    InMux I__2813 (
            .O(N__18623),
            .I(N__18594));
    InMux I__2812 (
            .O(N__18622),
            .I(N__18594));
    Span4Mux_v I__2811 (
            .O(N__18619),
            .I(N__18585));
    LocalMux I__2810 (
            .O(N__18616),
            .I(N__18585));
    Span4Mux_v I__2809 (
            .O(N__18613),
            .I(N__18585));
    Span4Mux_v I__2808 (
            .O(N__18608),
            .I(N__18585));
    InMux I__2807 (
            .O(N__18607),
            .I(N__18582));
    Odrv12 I__2806 (
            .O(N__18604),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2805 (
            .O(N__18599),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2804 (
            .O(N__18594),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__2803 (
            .O(N__18585),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    LocalMux I__2802 (
            .O(N__18582),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__2801 (
            .O(N__18571),
            .I(N__18567));
    InMux I__2800 (
            .O(N__18570),
            .I(N__18564));
    LocalMux I__2799 (
            .O(N__18567),
            .I(N__18560));
    LocalMux I__2798 (
            .O(N__18564),
            .I(N__18557));
    InMux I__2797 (
            .O(N__18563),
            .I(N__18554));
    Odrv4 I__2796 (
            .O(N__18560),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    Odrv4 I__2795 (
            .O(N__18557),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    LocalMux I__2794 (
            .O(N__18554),
            .I(\this_vga_signals.mult1_un68_sum_axbxc1 ));
    CascadeMux I__2793 (
            .O(N__18547),
            .I(N__18543));
    CascadeMux I__2792 (
            .O(N__18546),
            .I(N__18539));
    InMux I__2791 (
            .O(N__18543),
            .I(N__18536));
    InMux I__2790 (
            .O(N__18542),
            .I(N__18529));
    InMux I__2789 (
            .O(N__18539),
            .I(N__18529));
    LocalMux I__2788 (
            .O(N__18536),
            .I(N__18520));
    InMux I__2787 (
            .O(N__18535),
            .I(N__18517));
    InMux I__2786 (
            .O(N__18534),
            .I(N__18514));
    LocalMux I__2785 (
            .O(N__18529),
            .I(N__18511));
    CascadeMux I__2784 (
            .O(N__18528),
            .I(N__18508));
    CascadeMux I__2783 (
            .O(N__18527),
            .I(N__18504));
    CascadeMux I__2782 (
            .O(N__18526),
            .I(N__18501));
    CascadeMux I__2781 (
            .O(N__18525),
            .I(N__18497));
    CascadeMux I__2780 (
            .O(N__18524),
            .I(N__18494));
    InMux I__2779 (
            .O(N__18523),
            .I(N__18491));
    Span12Mux_h I__2778 (
            .O(N__18520),
            .I(N__18488));
    LocalMux I__2777 (
            .O(N__18517),
            .I(N__18481));
    LocalMux I__2776 (
            .O(N__18514),
            .I(N__18481));
    Span4Mux_h I__2775 (
            .O(N__18511),
            .I(N__18481));
    InMux I__2774 (
            .O(N__18508),
            .I(N__18478));
    InMux I__2773 (
            .O(N__18507),
            .I(N__18473));
    InMux I__2772 (
            .O(N__18504),
            .I(N__18473));
    InMux I__2771 (
            .O(N__18501),
            .I(N__18470));
    InMux I__2770 (
            .O(N__18500),
            .I(N__18463));
    InMux I__2769 (
            .O(N__18497),
            .I(N__18463));
    InMux I__2768 (
            .O(N__18494),
            .I(N__18463));
    LocalMux I__2767 (
            .O(N__18491),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv12 I__2766 (
            .O(N__18488),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__2765 (
            .O(N__18481),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2764 (
            .O(N__18478),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2763 (
            .O(N__18473),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2762 (
            .O(N__18470),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    LocalMux I__2761 (
            .O(N__18463),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__2760 (
            .O(N__18448),
            .I(N__18445));
    LocalMux I__2759 (
            .O(N__18445),
            .I(N__18438));
    InMux I__2758 (
            .O(N__18444),
            .I(N__18435));
    InMux I__2757 (
            .O(N__18443),
            .I(N__18430));
    InMux I__2756 (
            .O(N__18442),
            .I(N__18430));
    InMux I__2755 (
            .O(N__18441),
            .I(N__18424));
    Span4Mux_v I__2754 (
            .O(N__18438),
            .I(N__18417));
    LocalMux I__2753 (
            .O(N__18435),
            .I(N__18417));
    LocalMux I__2752 (
            .O(N__18430),
            .I(N__18417));
    InMux I__2751 (
            .O(N__18429),
            .I(N__18412));
    InMux I__2750 (
            .O(N__18428),
            .I(N__18412));
    InMux I__2749 (
            .O(N__18427),
            .I(N__18409));
    LocalMux I__2748 (
            .O(N__18424),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    Odrv4 I__2747 (
            .O(N__18417),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__2746 (
            .O(N__18412),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    LocalMux I__2745 (
            .O(N__18409),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3 ));
    InMux I__2744 (
            .O(N__18400),
            .I(N__18394));
    InMux I__2743 (
            .O(N__18399),
            .I(N__18390));
    InMux I__2742 (
            .O(N__18398),
            .I(N__18385));
    InMux I__2741 (
            .O(N__18397),
            .I(N__18385));
    LocalMux I__2740 (
            .O(N__18394),
            .I(N__18380));
    InMux I__2739 (
            .O(N__18393),
            .I(N__18377));
    LocalMux I__2738 (
            .O(N__18390),
            .I(N__18370));
    LocalMux I__2737 (
            .O(N__18385),
            .I(N__18370));
    InMux I__2736 (
            .O(N__18384),
            .I(N__18365));
    InMux I__2735 (
            .O(N__18383),
            .I(N__18365));
    Span4Mux_h I__2734 (
            .O(N__18380),
            .I(N__18359));
    LocalMux I__2733 (
            .O(N__18377),
            .I(N__18359));
    InMux I__2732 (
            .O(N__18376),
            .I(N__18356));
    InMux I__2731 (
            .O(N__18375),
            .I(N__18353));
    Span4Mux_v I__2730 (
            .O(N__18370),
            .I(N__18348));
    LocalMux I__2729 (
            .O(N__18365),
            .I(N__18348));
    InMux I__2728 (
            .O(N__18364),
            .I(N__18345));
    Odrv4 I__2727 (
            .O(N__18359),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2726 (
            .O(N__18356),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2725 (
            .O(N__18353),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv4 I__2724 (
            .O(N__18348),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__2723 (
            .O(N__18345),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    CascadeMux I__2722 (
            .O(N__18334),
            .I(\this_vga_signals.if_N_8_i_cascade_ ));
    InMux I__2721 (
            .O(N__18331),
            .I(N__18326));
    InMux I__2720 (
            .O(N__18330),
            .I(N__18321));
    CascadeMux I__2719 (
            .O(N__18329),
            .I(N__18318));
    LocalMux I__2718 (
            .O(N__18326),
            .I(N__18314));
    InMux I__2717 (
            .O(N__18325),
            .I(N__18309));
    InMux I__2716 (
            .O(N__18324),
            .I(N__18309));
    LocalMux I__2715 (
            .O(N__18321),
            .I(N__18306));
    InMux I__2714 (
            .O(N__18318),
            .I(N__18301));
    InMux I__2713 (
            .O(N__18317),
            .I(N__18301));
    Odrv4 I__2712 (
            .O(N__18314),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2711 (
            .O(N__18309),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv12 I__2710 (
            .O(N__18306),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__2709 (
            .O(N__18301),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    InMux I__2708 (
            .O(N__18292),
            .I(N__18289));
    LocalMux I__2707 (
            .O(N__18289),
            .I(\this_vga_signals.if_N_9_1 ));
    CascadeMux I__2706 (
            .O(N__18286),
            .I(\this_vga_signals.M_pcounter_q_3_1_cascade_ ));
    InMux I__2705 (
            .O(N__18283),
            .I(N__18278));
    InMux I__2704 (
            .O(N__18282),
            .I(N__18273));
    InMux I__2703 (
            .O(N__18281),
            .I(N__18273));
    LocalMux I__2702 (
            .O(N__18278),
            .I(\this_vga_signals.N_3_0 ));
    LocalMux I__2701 (
            .O(N__18273),
            .I(\this_vga_signals.N_3_0 ));
    InMux I__2700 (
            .O(N__18268),
            .I(N__18264));
    InMux I__2699 (
            .O(N__18267),
            .I(N__18261));
    LocalMux I__2698 (
            .O(N__18264),
            .I(N__18255));
    LocalMux I__2697 (
            .O(N__18261),
            .I(N__18255));
    CascadeMux I__2696 (
            .O(N__18260),
            .I(N__18252));
    Span4Mux_v I__2695 (
            .O(N__18255),
            .I(N__18248));
    InMux I__2694 (
            .O(N__18252),
            .I(N__18243));
    InMux I__2693 (
            .O(N__18251),
            .I(N__18243));
    Odrv4 I__2692 (
            .O(N__18248),
            .I(\this_vga_signals.SUM_3_i_0_0 ));
    LocalMux I__2691 (
            .O(N__18243),
            .I(\this_vga_signals.SUM_3_i_0_0 ));
    InMux I__2690 (
            .O(N__18238),
            .I(N__18235));
    LocalMux I__2689 (
            .O(N__18235),
            .I(N__18230));
    InMux I__2688 (
            .O(N__18234),
            .I(N__18225));
    InMux I__2687 (
            .O(N__18233),
            .I(N__18225));
    Odrv4 I__2686 (
            .O(N__18230),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ));
    LocalMux I__2685 (
            .O(N__18225),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ));
    InMux I__2684 (
            .O(N__18220),
            .I(N__18217));
    LocalMux I__2683 (
            .O(N__18217),
            .I(N__18214));
    Odrv12 I__2682 (
            .O(N__18214),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0 ));
    CascadeMux I__2681 (
            .O(N__18211),
            .I(N__18205));
    InMux I__2680 (
            .O(N__18210),
            .I(N__18201));
    InMux I__2679 (
            .O(N__18209),
            .I(N__18198));
    InMux I__2678 (
            .O(N__18208),
            .I(N__18191));
    InMux I__2677 (
            .O(N__18205),
            .I(N__18191));
    CascadeMux I__2676 (
            .O(N__18204),
            .I(N__18188));
    LocalMux I__2675 (
            .O(N__18201),
            .I(N__18182));
    LocalMux I__2674 (
            .O(N__18198),
            .I(N__18179));
    InMux I__2673 (
            .O(N__18197),
            .I(N__18176));
    InMux I__2672 (
            .O(N__18196),
            .I(N__18173));
    LocalMux I__2671 (
            .O(N__18191),
            .I(N__18170));
    InMux I__2670 (
            .O(N__18188),
            .I(N__18167));
    InMux I__2669 (
            .O(N__18187),
            .I(N__18160));
    InMux I__2668 (
            .O(N__18186),
            .I(N__18160));
    InMux I__2667 (
            .O(N__18185),
            .I(N__18160));
    Odrv4 I__2666 (
            .O(N__18182),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2665 (
            .O(N__18179),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2664 (
            .O(N__18176),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2663 (
            .O(N__18173),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__2662 (
            .O(N__18170),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2661 (
            .O(N__18167),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__2660 (
            .O(N__18160),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__2659 (
            .O(N__18145),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ));
    InMux I__2658 (
            .O(N__18142),
            .I(N__18137));
    InMux I__2657 (
            .O(N__18141),
            .I(N__18134));
    InMux I__2656 (
            .O(N__18140),
            .I(N__18130));
    LocalMux I__2655 (
            .O(N__18137),
            .I(N__18124));
    LocalMux I__2654 (
            .O(N__18134),
            .I(N__18121));
    InMux I__2653 (
            .O(N__18133),
            .I(N__18118));
    LocalMux I__2652 (
            .O(N__18130),
            .I(N__18109));
    InMux I__2651 (
            .O(N__18129),
            .I(N__18106));
    InMux I__2650 (
            .O(N__18128),
            .I(N__18103));
    InMux I__2649 (
            .O(N__18127),
            .I(N__18100));
    Span4Mux_v I__2648 (
            .O(N__18124),
            .I(N__18093));
    Span4Mux_v I__2647 (
            .O(N__18121),
            .I(N__18093));
    LocalMux I__2646 (
            .O(N__18118),
            .I(N__18093));
    InMux I__2645 (
            .O(N__18117),
            .I(N__18086));
    InMux I__2644 (
            .O(N__18116),
            .I(N__18086));
    InMux I__2643 (
            .O(N__18115),
            .I(N__18086));
    InMux I__2642 (
            .O(N__18114),
            .I(N__18079));
    InMux I__2641 (
            .O(N__18113),
            .I(N__18079));
    InMux I__2640 (
            .O(N__18112),
            .I(N__18079));
    Odrv12 I__2639 (
            .O(N__18109),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2638 (
            .O(N__18106),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2637 (
            .O(N__18103),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2636 (
            .O(N__18100),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__2635 (
            .O(N__18093),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2634 (
            .O(N__18086),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__2633 (
            .O(N__18079),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__2632 (
            .O(N__18064),
            .I(N__18061));
    LocalMux I__2631 (
            .O(N__18061),
            .I(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ));
    CascadeMux I__2630 (
            .O(N__18058),
            .I(N__18053));
    InMux I__2629 (
            .O(N__18057),
            .I(N__18040));
    InMux I__2628 (
            .O(N__18056),
            .I(N__18040));
    InMux I__2627 (
            .O(N__18053),
            .I(N__18040));
    InMux I__2626 (
            .O(N__18052),
            .I(N__18040));
    InMux I__2625 (
            .O(N__18051),
            .I(N__18037));
    InMux I__2624 (
            .O(N__18050),
            .I(N__18034));
    InMux I__2623 (
            .O(N__18049),
            .I(N__18031));
    LocalMux I__2622 (
            .O(N__18040),
            .I(N__18024));
    LocalMux I__2621 (
            .O(N__18037),
            .I(N__18024));
    LocalMux I__2620 (
            .O(N__18034),
            .I(N__18024));
    LocalMux I__2619 (
            .O(N__18031),
            .I(N_28_0));
    Odrv12 I__2618 (
            .O(N__18024),
            .I(N_28_0));
    InMux I__2617 (
            .O(N__18019),
            .I(N__18016));
    LocalMux I__2616 (
            .O(N__18016),
            .I(\this_vga_signals.M_hcounter_d7lt7_0 ));
    CascadeMux I__2615 (
            .O(N__18013),
            .I(N__18010));
    InMux I__2614 (
            .O(N__18010),
            .I(N__18007));
    LocalMux I__2613 (
            .O(N__18007),
            .I(N__18004));
    Span4Mux_s2_v I__2612 (
            .O(N__18004),
            .I(N__18001));
    Odrv4 I__2611 (
            .O(N__18001),
            .I(M_this_vga_signals_address_5));
    InMux I__2610 (
            .O(N__17998),
            .I(N__17987));
    InMux I__2609 (
            .O(N__17997),
            .I(N__17987));
    InMux I__2608 (
            .O(N__17996),
            .I(N__17987));
    InMux I__2607 (
            .O(N__17995),
            .I(N__17984));
    InMux I__2606 (
            .O(N__17994),
            .I(N__17981));
    LocalMux I__2605 (
            .O(N__17987),
            .I(N__17978));
    LocalMux I__2604 (
            .O(N__17984),
            .I(N__17973));
    LocalMux I__2603 (
            .O(N__17981),
            .I(N__17973));
    Span4Mux_h I__2602 (
            .O(N__17978),
            .I(N__17970));
    Span4Mux_h I__2601 (
            .O(N__17973),
            .I(N__17967));
    Odrv4 I__2600 (
            .O(N__17970),
            .I(M_this_vram_read_data_2));
    Odrv4 I__2599 (
            .O(N__17967),
            .I(M_this_vram_read_data_2));
    CascadeMux I__2598 (
            .O(N__17962),
            .I(N__17957));
    CascadeMux I__2597 (
            .O(N__17961),
            .I(N__17953));
    InMux I__2596 (
            .O(N__17960),
            .I(N__17949));
    InMux I__2595 (
            .O(N__17957),
            .I(N__17944));
    InMux I__2594 (
            .O(N__17956),
            .I(N__17944));
    InMux I__2593 (
            .O(N__17953),
            .I(N__17940));
    InMux I__2592 (
            .O(N__17952),
            .I(N__17937));
    LocalMux I__2591 (
            .O(N__17949),
            .I(N__17934));
    LocalMux I__2590 (
            .O(N__17944),
            .I(N__17931));
    InMux I__2589 (
            .O(N__17943),
            .I(N__17928));
    LocalMux I__2588 (
            .O(N__17940),
            .I(N__17925));
    LocalMux I__2587 (
            .O(N__17937),
            .I(N__17922));
    Span4Mux_h I__2586 (
            .O(N__17934),
            .I(N__17919));
    Span4Mux_h I__2585 (
            .O(N__17931),
            .I(N__17912));
    LocalMux I__2584 (
            .O(N__17928),
            .I(N__17912));
    Span4Mux_h I__2583 (
            .O(N__17925),
            .I(N__17912));
    Span4Mux_h I__2582 (
            .O(N__17922),
            .I(N__17909));
    Odrv4 I__2581 (
            .O(N__17919),
            .I(M_this_vram_read_data_1));
    Odrv4 I__2580 (
            .O(N__17912),
            .I(M_this_vram_read_data_1));
    Odrv4 I__2579 (
            .O(N__17909),
            .I(M_this_vram_read_data_1));
    CascadeMux I__2578 (
            .O(N__17902),
            .I(N__17898));
    CascadeMux I__2577 (
            .O(N__17901),
            .I(N__17894));
    InMux I__2576 (
            .O(N__17898),
            .I(N__17888));
    InMux I__2575 (
            .O(N__17897),
            .I(N__17885));
    InMux I__2574 (
            .O(N__17894),
            .I(N__17882));
    InMux I__2573 (
            .O(N__17893),
            .I(N__17875));
    InMux I__2572 (
            .O(N__17892),
            .I(N__17875));
    InMux I__2571 (
            .O(N__17891),
            .I(N__17875));
    LocalMux I__2570 (
            .O(N__17888),
            .I(N__17866));
    LocalMux I__2569 (
            .O(N__17885),
            .I(N__17866));
    LocalMux I__2568 (
            .O(N__17882),
            .I(N__17866));
    LocalMux I__2567 (
            .O(N__17875),
            .I(N__17866));
    Span4Mux_v I__2566 (
            .O(N__17866),
            .I(N__17863));
    Span4Mux_h I__2565 (
            .O(N__17863),
            .I(N__17860));
    Odrv4 I__2564 (
            .O(N__17860),
            .I(M_this_vram_read_data_0));
    CascadeMux I__2563 (
            .O(N__17857),
            .I(N__17854));
    InMux I__2562 (
            .O(N__17854),
            .I(N__17847));
    InMux I__2561 (
            .O(N__17853),
            .I(N__17847));
    CascadeMux I__2560 (
            .O(N__17852),
            .I(N__17843));
    LocalMux I__2559 (
            .O(N__17847),
            .I(N__17838));
    InMux I__2558 (
            .O(N__17846),
            .I(N__17835));
    InMux I__2557 (
            .O(N__17843),
            .I(N__17832));
    InMux I__2556 (
            .O(N__17842),
            .I(N__17829));
    InMux I__2555 (
            .O(N__17841),
            .I(N__17826));
    Span4Mux_v I__2554 (
            .O(N__17838),
            .I(N__17823));
    LocalMux I__2553 (
            .O(N__17835),
            .I(N__17814));
    LocalMux I__2552 (
            .O(N__17832),
            .I(N__17814));
    LocalMux I__2551 (
            .O(N__17829),
            .I(N__17814));
    LocalMux I__2550 (
            .O(N__17826),
            .I(N__17814));
    Span4Mux_h I__2549 (
            .O(N__17823),
            .I(N__17809));
    Span4Mux_v I__2548 (
            .O(N__17814),
            .I(N__17809));
    Sp12to4 I__2547 (
            .O(N__17809),
            .I(N__17806));
    Odrv12 I__2546 (
            .O(N__17806),
            .I(M_this_vram_read_data_3));
    InMux I__2545 (
            .O(N__17803),
            .I(N__17800));
    LocalMux I__2544 (
            .O(N__17800),
            .I(N__17797));
    Span4Mux_v I__2543 (
            .O(N__17797),
            .I(N__17794));
    Odrv4 I__2542 (
            .O(N__17794),
            .I(\this_vga_ramdac.i2_mux_0 ));
    CascadeMux I__2541 (
            .O(N__17791),
            .I(\this_vga_signals.N_2_8_0_cascade_ ));
    InMux I__2540 (
            .O(N__17788),
            .I(N__17785));
    LocalMux I__2539 (
            .O(N__17785),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_2_am ));
    InMux I__2538 (
            .O(N__17782),
            .I(N__17779));
    LocalMux I__2537 (
            .O(N__17779),
            .I(N__17776));
    Odrv4 I__2536 (
            .O(N__17776),
            .I(\this_vga_signals.haddress_1Z0Z_0 ));
    InMux I__2535 (
            .O(N__17773),
            .I(N__17767));
    InMux I__2534 (
            .O(N__17772),
            .I(N__17767));
    LocalMux I__2533 (
            .O(N__17767),
            .I(N__17762));
    InMux I__2532 (
            .O(N__17766),
            .I(N__17757));
    InMux I__2531 (
            .O(N__17765),
            .I(N__17757));
    Odrv4 I__2530 (
            .O(N__17762),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__2529 (
            .O(N__17757),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    InMux I__2528 (
            .O(N__17752),
            .I(N__17749));
    LocalMux I__2527 (
            .O(N__17749),
            .I(N__17746));
    Odrv4 I__2526 (
            .O(N__17746),
            .I(\this_vga_signals.mult1_un89_sum_c3 ));
    CascadeMux I__2525 (
            .O(N__17743),
            .I(N__17740));
    InMux I__2524 (
            .O(N__17740),
            .I(N__17734));
    InMux I__2523 (
            .O(N__17739),
            .I(N__17734));
    LocalMux I__2522 (
            .O(N__17734),
            .I(N__17730));
    InMux I__2521 (
            .O(N__17733),
            .I(N__17727));
    Span4Mux_h I__2520 (
            .O(N__17730),
            .I(N__17724));
    LocalMux I__2519 (
            .O(N__17727),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    Odrv4 I__2518 (
            .O(N__17724),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_0 ));
    InMux I__2517 (
            .O(N__17719),
            .I(N__17716));
    LocalMux I__2516 (
            .O(N__17716),
            .I(N__17712));
    InMux I__2515 (
            .O(N__17715),
            .I(N__17709));
    Span4Mux_v I__2514 (
            .O(N__17712),
            .I(N__17699));
    LocalMux I__2513 (
            .O(N__17709),
            .I(N__17699));
    InMux I__2512 (
            .O(N__17708),
            .I(N__17692));
    InMux I__2511 (
            .O(N__17707),
            .I(N__17692));
    InMux I__2510 (
            .O(N__17706),
            .I(N__17692));
    InMux I__2509 (
            .O(N__17705),
            .I(N__17687));
    InMux I__2508 (
            .O(N__17704),
            .I(N__17687));
    Span4Mux_v I__2507 (
            .O(N__17699),
            .I(N__17682));
    LocalMux I__2506 (
            .O(N__17692),
            .I(N__17682));
    LocalMux I__2505 (
            .O(N__17687),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    Odrv4 I__2504 (
            .O(N__17682),
            .I(\this_vga_signals.mult1_un61_sum_0_3 ));
    InMux I__2503 (
            .O(N__17677),
            .I(N__17674));
    LocalMux I__2502 (
            .O(N__17674),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_2_bm ));
    InMux I__2501 (
            .O(N__17671),
            .I(N__17667));
    InMux I__2500 (
            .O(N__17670),
            .I(N__17664));
    LocalMux I__2499 (
            .O(N__17667),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    LocalMux I__2498 (
            .O(N__17664),
            .I(\this_vga_signals.mult1_un75_sum_c2_0 ));
    InMux I__2497 (
            .O(N__17659),
            .I(N__17656));
    LocalMux I__2496 (
            .O(N__17656),
            .I(N__17653));
    Odrv4 I__2495 (
            .O(N__17653),
            .I(\this_vga_ramdac.i2_mux ));
    InMux I__2494 (
            .O(N__17650),
            .I(N__17647));
    LocalMux I__2493 (
            .O(N__17647),
            .I(N__17639));
    InMux I__2492 (
            .O(N__17646),
            .I(N__17634));
    InMux I__2491 (
            .O(N__17645),
            .I(N__17634));
    InMux I__2490 (
            .O(N__17644),
            .I(N__17627));
    InMux I__2489 (
            .O(N__17643),
            .I(N__17627));
    InMux I__2488 (
            .O(N__17642),
            .I(N__17627));
    Odrv4 I__2487 (
            .O(N__17639),
            .I(M_pcounter_q_ret_1_RNI4VLK7));
    LocalMux I__2486 (
            .O(N__17634),
            .I(M_pcounter_q_ret_1_RNI4VLK7));
    LocalMux I__2485 (
            .O(N__17627),
            .I(M_pcounter_q_ret_1_RNI4VLK7));
    InMux I__2484 (
            .O(N__17620),
            .I(N__17617));
    LocalMux I__2483 (
            .O(N__17617),
            .I(N__17613));
    CascadeMux I__2482 (
            .O(N__17616),
            .I(N__17610));
    Span12Mux_v I__2481 (
            .O(N__17613),
            .I(N__17607));
    InMux I__2480 (
            .O(N__17610),
            .I(N__17604));
    Odrv12 I__2479 (
            .O(N__17607),
            .I(\this_vga_ramdac.N_2688_reto ));
    LocalMux I__2478 (
            .O(N__17604),
            .I(\this_vga_ramdac.N_2688_reto ));
    InMux I__2477 (
            .O(N__17599),
            .I(N__17591));
    CascadeMux I__2476 (
            .O(N__17598),
            .I(N__17587));
    CascadeMux I__2475 (
            .O(N__17597),
            .I(N__17580));
    InMux I__2474 (
            .O(N__17596),
            .I(N__17577));
    InMux I__2473 (
            .O(N__17595),
            .I(N__17573));
    InMux I__2472 (
            .O(N__17594),
            .I(N__17560));
    LocalMux I__2471 (
            .O(N__17591),
            .I(N__17557));
    InMux I__2470 (
            .O(N__17590),
            .I(N__17554));
    InMux I__2469 (
            .O(N__17587),
            .I(N__17551));
    InMux I__2468 (
            .O(N__17586),
            .I(N__17546));
    InMux I__2467 (
            .O(N__17585),
            .I(N__17546));
    InMux I__2466 (
            .O(N__17584),
            .I(N__17543));
    InMux I__2465 (
            .O(N__17583),
            .I(N__17540));
    InMux I__2464 (
            .O(N__17580),
            .I(N__17537));
    LocalMux I__2463 (
            .O(N__17577),
            .I(N__17534));
    CascadeMux I__2462 (
            .O(N__17576),
            .I(N__17531));
    LocalMux I__2461 (
            .O(N__17573),
            .I(N__17526));
    InMux I__2460 (
            .O(N__17572),
            .I(N__17521));
    InMux I__2459 (
            .O(N__17571),
            .I(N__17521));
    InMux I__2458 (
            .O(N__17570),
            .I(N__17517));
    CascadeMux I__2457 (
            .O(N__17569),
            .I(N__17513));
    InMux I__2456 (
            .O(N__17568),
            .I(N__17503));
    InMux I__2455 (
            .O(N__17567),
            .I(N__17503));
    InMux I__2454 (
            .O(N__17566),
            .I(N__17503));
    InMux I__2453 (
            .O(N__17565),
            .I(N__17503));
    InMux I__2452 (
            .O(N__17564),
            .I(N__17498));
    InMux I__2451 (
            .O(N__17563),
            .I(N__17498));
    LocalMux I__2450 (
            .O(N__17560),
            .I(N__17495));
    Span4Mux_h I__2449 (
            .O(N__17557),
            .I(N__17492));
    LocalMux I__2448 (
            .O(N__17554),
            .I(N__17485));
    LocalMux I__2447 (
            .O(N__17551),
            .I(N__17485));
    LocalMux I__2446 (
            .O(N__17546),
            .I(N__17485));
    LocalMux I__2445 (
            .O(N__17543),
            .I(N__17482));
    LocalMux I__2444 (
            .O(N__17540),
            .I(N__17479));
    LocalMux I__2443 (
            .O(N__17537),
            .I(N__17476));
    Span4Mux_v I__2442 (
            .O(N__17534),
            .I(N__17472));
    InMux I__2441 (
            .O(N__17531),
            .I(N__17467));
    InMux I__2440 (
            .O(N__17530),
            .I(N__17467));
    InMux I__2439 (
            .O(N__17529),
            .I(N__17464));
    Span4Mux_v I__2438 (
            .O(N__17526),
            .I(N__17459));
    LocalMux I__2437 (
            .O(N__17521),
            .I(N__17459));
    InMux I__2436 (
            .O(N__17520),
            .I(N__17456));
    LocalMux I__2435 (
            .O(N__17517),
            .I(N__17453));
    InMux I__2434 (
            .O(N__17516),
            .I(N__17446));
    InMux I__2433 (
            .O(N__17513),
            .I(N__17446));
    InMux I__2432 (
            .O(N__17512),
            .I(N__17446));
    LocalMux I__2431 (
            .O(N__17503),
            .I(N__17437));
    LocalMux I__2430 (
            .O(N__17498),
            .I(N__17437));
    Span4Mux_h I__2429 (
            .O(N__17495),
            .I(N__17437));
    Span4Mux_h I__2428 (
            .O(N__17492),
            .I(N__17437));
    Span4Mux_v I__2427 (
            .O(N__17485),
            .I(N__17428));
    Span4Mux_h I__2426 (
            .O(N__17482),
            .I(N__17428));
    Span4Mux_v I__2425 (
            .O(N__17479),
            .I(N__17428));
    Span4Mux_v I__2424 (
            .O(N__17476),
            .I(N__17428));
    InMux I__2423 (
            .O(N__17475),
            .I(N__17425));
    Odrv4 I__2422 (
            .O(N__17472),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2421 (
            .O(N__17467),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2420 (
            .O(N__17464),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2419 (
            .O(N__17459),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2418 (
            .O(N__17456),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2417 (
            .O(N__17453),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2416 (
            .O(N__17446),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2415 (
            .O(N__17437),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__2414 (
            .O(N__17428),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__2413 (
            .O(N__17425),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    InMux I__2412 (
            .O(N__17404),
            .I(N__17400));
    CascadeMux I__2411 (
            .O(N__17403),
            .I(N__17396));
    LocalMux I__2410 (
            .O(N__17400),
            .I(N__17386));
    InMux I__2409 (
            .O(N__17399),
            .I(N__17381));
    InMux I__2408 (
            .O(N__17396),
            .I(N__17381));
    CascadeMux I__2407 (
            .O(N__17395),
            .I(N__17376));
    InMux I__2406 (
            .O(N__17394),
            .I(N__17372));
    InMux I__2405 (
            .O(N__17393),
            .I(N__17369));
    InMux I__2404 (
            .O(N__17392),
            .I(N__17365));
    InMux I__2403 (
            .O(N__17391),
            .I(N__17362));
    InMux I__2402 (
            .O(N__17390),
            .I(N__17359));
    InMux I__2401 (
            .O(N__17389),
            .I(N__17356));
    Span4Mux_v I__2400 (
            .O(N__17386),
            .I(N__17351));
    LocalMux I__2399 (
            .O(N__17381),
            .I(N__17351));
    CascadeMux I__2398 (
            .O(N__17380),
            .I(N__17347));
    InMux I__2397 (
            .O(N__17379),
            .I(N__17340));
    InMux I__2396 (
            .O(N__17376),
            .I(N__17335));
    InMux I__2395 (
            .O(N__17375),
            .I(N__17335));
    LocalMux I__2394 (
            .O(N__17372),
            .I(N__17330));
    LocalMux I__2393 (
            .O(N__17369),
            .I(N__17330));
    InMux I__2392 (
            .O(N__17368),
            .I(N__17327));
    LocalMux I__2391 (
            .O(N__17365),
            .I(N__17322));
    LocalMux I__2390 (
            .O(N__17362),
            .I(N__17319));
    LocalMux I__2389 (
            .O(N__17359),
            .I(N__17314));
    LocalMux I__2388 (
            .O(N__17356),
            .I(N__17314));
    Span4Mux_v I__2387 (
            .O(N__17351),
            .I(N__17311));
    InMux I__2386 (
            .O(N__17350),
            .I(N__17306));
    InMux I__2385 (
            .O(N__17347),
            .I(N__17306));
    InMux I__2384 (
            .O(N__17346),
            .I(N__17301));
    InMux I__2383 (
            .O(N__17345),
            .I(N__17301));
    InMux I__2382 (
            .O(N__17344),
            .I(N__17298));
    InMux I__2381 (
            .O(N__17343),
            .I(N__17295));
    LocalMux I__2380 (
            .O(N__17340),
            .I(N__17292));
    LocalMux I__2379 (
            .O(N__17335),
            .I(N__17289));
    Span4Mux_v I__2378 (
            .O(N__17330),
            .I(N__17284));
    LocalMux I__2377 (
            .O(N__17327),
            .I(N__17284));
    InMux I__2376 (
            .O(N__17326),
            .I(N__17279));
    InMux I__2375 (
            .O(N__17325),
            .I(N__17279));
    Span4Mux_s1_h I__2374 (
            .O(N__17322),
            .I(N__17270));
    Span4Mux_v I__2373 (
            .O(N__17319),
            .I(N__17270));
    Span4Mux_v I__2372 (
            .O(N__17314),
            .I(N__17270));
    Span4Mux_s1_h I__2371 (
            .O(N__17311),
            .I(N__17270));
    LocalMux I__2370 (
            .O(N__17306),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2369 (
            .O(N__17301),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2368 (
            .O(N__17298),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2367 (
            .O(N__17295),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2366 (
            .O(N__17292),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2365 (
            .O(N__17289),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2364 (
            .O(N__17284),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    LocalMux I__2363 (
            .O(N__17279),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    Odrv4 I__2362 (
            .O(N__17270),
            .I(\this_vga_signals.M_vcounter_qZ0Z_6 ));
    CascadeMux I__2361 (
            .O(N__17251),
            .I(N__17248));
    InMux I__2360 (
            .O(N__17248),
            .I(N__17245));
    LocalMux I__2359 (
            .O(N__17245),
            .I(N__17242));
    Span4Mux_h I__2358 (
            .O(N__17242),
            .I(N__17239));
    Odrv4 I__2357 (
            .O(N__17239),
            .I(\this_vga_signals.g0_6_0_0 ));
    IoInMux I__2356 (
            .O(N__17236),
            .I(N__17233));
    LocalMux I__2355 (
            .O(N__17233),
            .I(N__17230));
    Span4Mux_s3_v I__2354 (
            .O(N__17230),
            .I(N__17227));
    Span4Mux_v I__2353 (
            .O(N__17227),
            .I(N__17224));
    Sp12to4 I__2352 (
            .O(N__17224),
            .I(N__17221));
    Span12Mux_s5_h I__2351 (
            .O(N__17221),
            .I(N__17218));
    Odrv12 I__2350 (
            .O(N__17218),
            .I(M_hcounter_q_esr_RNIU8TO_9));
    CascadeMux I__2349 (
            .O(N__17215),
            .I(N__17212));
    InMux I__2348 (
            .O(N__17212),
            .I(N__17209));
    LocalMux I__2347 (
            .O(N__17209),
            .I(M_this_vga_signals_address_2));
    CascadeMux I__2346 (
            .O(N__17206),
            .I(N__17203));
    InMux I__2345 (
            .O(N__17203),
            .I(N__17200));
    LocalMux I__2344 (
            .O(N__17200),
            .I(M_this_vga_signals_address_0));
    CascadeMux I__2343 (
            .O(N__17197),
            .I(N__17194));
    InMux I__2342 (
            .O(N__17194),
            .I(N__17191));
    LocalMux I__2341 (
            .O(N__17191),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__2340 (
            .O(N__17188),
            .I(N__17185));
    InMux I__2339 (
            .O(N__17185),
            .I(N__17182));
    LocalMux I__2338 (
            .O(N__17182),
            .I(M_this_vga_signals_address_4));
    InMux I__2337 (
            .O(N__17179),
            .I(N__17173));
    InMux I__2336 (
            .O(N__17178),
            .I(N__17173));
    LocalMux I__2335 (
            .O(N__17173),
            .I(N__17170));
    Span4Mux_h I__2334 (
            .O(N__17170),
            .I(N__17167));
    Odrv4 I__2333 (
            .O(N__17167),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ));
    CascadeMux I__2332 (
            .O(N__17164),
            .I(N__17161));
    InMux I__2331 (
            .O(N__17161),
            .I(N__17158));
    LocalMux I__2330 (
            .O(N__17158),
            .I(N__17155));
    Odrv4 I__2329 (
            .O(N__17155),
            .I(M_this_vga_signals_address_1));
    InMux I__2328 (
            .O(N__17152),
            .I(N__17149));
    LocalMux I__2327 (
            .O(N__17149),
            .I(\this_vga_signals.M_hcounter_d7lt4 ));
    InMux I__2326 (
            .O(N__17146),
            .I(N__17143));
    LocalMux I__2325 (
            .O(N__17143),
            .I(N__17140));
    Span4Mux_v I__2324 (
            .O(N__17140),
            .I(N__17136));
    CascadeMux I__2323 (
            .O(N__17139),
            .I(N__17133));
    Span4Mux_v I__2322 (
            .O(N__17136),
            .I(N__17130));
    InMux I__2321 (
            .O(N__17133),
            .I(N__17127));
    Odrv4 I__2320 (
            .O(N__17130),
            .I(\this_vga_ramdac.N_2691_reto ));
    LocalMux I__2319 (
            .O(N__17127),
            .I(\this_vga_ramdac.N_2691_reto ));
    InMux I__2318 (
            .O(N__17122),
            .I(N__17119));
    LocalMux I__2317 (
            .O(N__17119),
            .I(N__17116));
    Odrv4 I__2316 (
            .O(N__17116),
            .I(\this_vga_ramdac.m16 ));
    InMux I__2315 (
            .O(N__17113),
            .I(N__17110));
    LocalMux I__2314 (
            .O(N__17110),
            .I(N__17107));
    Span4Mux_h I__2313 (
            .O(N__17107),
            .I(N__17103));
    CascadeMux I__2312 (
            .O(N__17106),
            .I(N__17100));
    Span4Mux_v I__2311 (
            .O(N__17103),
            .I(N__17097));
    InMux I__2310 (
            .O(N__17100),
            .I(N__17094));
    Odrv4 I__2309 (
            .O(N__17097),
            .I(\this_vga_ramdac.N_2689_reto ));
    LocalMux I__2308 (
            .O(N__17094),
            .I(\this_vga_ramdac.N_2689_reto ));
    InMux I__2307 (
            .O(N__17089),
            .I(N__17086));
    LocalMux I__2306 (
            .O(N__17086),
            .I(N__17083));
    Odrv4 I__2305 (
            .O(N__17083),
            .I(\this_vga_signals.N_822_0 ));
    InMux I__2304 (
            .O(N__17080),
            .I(N__17077));
    LocalMux I__2303 (
            .O(N__17077),
            .I(N__17074));
    Odrv4 I__2302 (
            .O(N__17074),
            .I(\this_vga_signals.M_lcounter_q_3_i_o2_2_1_1 ));
    InMux I__2301 (
            .O(N__17071),
            .I(N__17068));
    LocalMux I__2300 (
            .O(N__17068),
            .I(N__17065));
    Odrv12 I__2299 (
            .O(N__17065),
            .I(\this_vga_ramdac.N_24_mux ));
    CascadeMux I__2298 (
            .O(N__17062),
            .I(M_pcounter_q_ret_1_RNI4VLK7_cascade_));
    InMux I__2297 (
            .O(N__17059),
            .I(N__17056));
    LocalMux I__2296 (
            .O(N__17056),
            .I(N__17053));
    Span4Mux_h I__2295 (
            .O(N__17053),
            .I(N__17049));
    InMux I__2294 (
            .O(N__17052),
            .I(N__17046));
    Odrv4 I__2293 (
            .O(N__17049),
            .I(\this_vga_ramdac.N_2686_reto ));
    LocalMux I__2292 (
            .O(N__17046),
            .I(\this_vga_ramdac.N_2686_reto ));
    CascadeMux I__2291 (
            .O(N__17041),
            .I(N__17038));
    InMux I__2290 (
            .O(N__17038),
            .I(N__17035));
    LocalMux I__2289 (
            .O(N__17035),
            .I(\this_vga_signals.mult1_un82_sum_c3 ));
    CascadeMux I__2288 (
            .O(N__17032),
            .I(\this_vga_signals.d_N_11_cascade_ ));
    InMux I__2287 (
            .O(N__17029),
            .I(N__17026));
    LocalMux I__2286 (
            .O(N__17026),
            .I(N__17023));
    Odrv4 I__2285 (
            .O(N__17023),
            .I(\this_vga_ramdac.m6 ));
    InMux I__2284 (
            .O(N__17020),
            .I(N__17016));
    CascadeMux I__2283 (
            .O(N__17019),
            .I(N__17013));
    LocalMux I__2282 (
            .O(N__17016),
            .I(N__17010));
    InMux I__2281 (
            .O(N__17013),
            .I(N__17007));
    Odrv12 I__2280 (
            .O(N__17010),
            .I(\this_vga_ramdac.N_2687_reto ));
    LocalMux I__2279 (
            .O(N__17007),
            .I(\this_vga_ramdac.N_2687_reto ));
    InMux I__2278 (
            .O(N__17002),
            .I(N__16998));
    InMux I__2277 (
            .O(N__17001),
            .I(N__16994));
    LocalMux I__2276 (
            .O(N__16998),
            .I(N__16989));
    InMux I__2275 (
            .O(N__16997),
            .I(N__16986));
    LocalMux I__2274 (
            .O(N__16994),
            .I(N__16983));
    InMux I__2273 (
            .O(N__16993),
            .I(N__16980));
    CascadeMux I__2272 (
            .O(N__16992),
            .I(N__16977));
    Span4Mux_v I__2271 (
            .O(N__16989),
            .I(N__16973));
    LocalMux I__2270 (
            .O(N__16986),
            .I(N__16970));
    Span4Mux_v I__2269 (
            .O(N__16983),
            .I(N__16965));
    LocalMux I__2268 (
            .O(N__16980),
            .I(N__16965));
    InMux I__2267 (
            .O(N__16977),
            .I(N__16960));
    InMux I__2266 (
            .O(N__16976),
            .I(N__16960));
    Span4Mux_h I__2265 (
            .O(N__16973),
            .I(N__16954));
    Span4Mux_v I__2264 (
            .O(N__16970),
            .I(N__16954));
    Span4Mux_v I__2263 (
            .O(N__16965),
            .I(N__16951));
    LocalMux I__2262 (
            .O(N__16960),
            .I(N__16948));
    CascadeMux I__2261 (
            .O(N__16959),
            .I(N__16945));
    Span4Mux_v I__2260 (
            .O(N__16954),
            .I(N__16942));
    Span4Mux_h I__2259 (
            .O(N__16951),
            .I(N__16939));
    Span12Mux_s8_v I__2258 (
            .O(N__16948),
            .I(N__16936));
    InMux I__2257 (
            .O(N__16945),
            .I(N__16933));
    Odrv4 I__2256 (
            .O(N__16942),
            .I(\this_vga_ramdac.N_28_i_reto ));
    Odrv4 I__2255 (
            .O(N__16939),
            .I(\this_vga_ramdac.N_28_i_reto ));
    Odrv12 I__2254 (
            .O(N__16936),
            .I(\this_vga_ramdac.N_28_i_reto ));
    LocalMux I__2253 (
            .O(N__16933),
            .I(\this_vga_ramdac.N_28_i_reto ));
    InMux I__2252 (
            .O(N__16924),
            .I(N__16921));
    LocalMux I__2251 (
            .O(N__16921),
            .I(N__16918));
    Odrv12 I__2250 (
            .O(N__16918),
            .I(\this_vga_ramdac.m19 ));
    InMux I__2249 (
            .O(N__16915),
            .I(N__16912));
    LocalMux I__2248 (
            .O(N__16912),
            .I(N__16909));
    Span4Mux_v I__2247 (
            .O(N__16909),
            .I(N__16905));
    CascadeMux I__2246 (
            .O(N__16908),
            .I(N__16902));
    Span4Mux_h I__2245 (
            .O(N__16905),
            .I(N__16899));
    InMux I__2244 (
            .O(N__16902),
            .I(N__16896));
    Odrv4 I__2243 (
            .O(N__16899),
            .I(\this_vga_ramdac.N_2690_reto ));
    LocalMux I__2242 (
            .O(N__16896),
            .I(\this_vga_ramdac.N_2690_reto ));
    InMux I__2241 (
            .O(N__16891),
            .I(N__16886));
    InMux I__2240 (
            .O(N__16890),
            .I(N__16881));
    InMux I__2239 (
            .O(N__16889),
            .I(N__16881));
    LocalMux I__2238 (
            .O(N__16886),
            .I(N__16878));
    LocalMux I__2237 (
            .O(N__16881),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    Odrv4 I__2236 (
            .O(N__16878),
            .I(\this_vga_signals.mult1_un61_sum_axb1 ));
    CascadeMux I__2235 (
            .O(N__16873),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ));
    CascadeMux I__2234 (
            .O(N__16870),
            .I(N__16866));
    InMux I__2233 (
            .O(N__16869),
            .I(N__16861));
    InMux I__2232 (
            .O(N__16866),
            .I(N__16861));
    LocalMux I__2231 (
            .O(N__16861),
            .I(N__16850));
    InMux I__2230 (
            .O(N__16860),
            .I(N__16847));
    CascadeMux I__2229 (
            .O(N__16859),
            .I(N__16843));
    CascadeMux I__2228 (
            .O(N__16858),
            .I(N__16837));
    InMux I__2227 (
            .O(N__16857),
            .I(N__16833));
    CascadeMux I__2226 (
            .O(N__16856),
            .I(N__16830));
    CascadeMux I__2225 (
            .O(N__16855),
            .I(N__16827));
    CascadeMux I__2224 (
            .O(N__16854),
            .I(N__16824));
    CascadeMux I__2223 (
            .O(N__16853),
            .I(N__16819));
    Span4Mux_v I__2222 (
            .O(N__16850),
            .I(N__16815));
    LocalMux I__2221 (
            .O(N__16847),
            .I(N__16812));
    InMux I__2220 (
            .O(N__16846),
            .I(N__16809));
    InMux I__2219 (
            .O(N__16843),
            .I(N__16804));
    InMux I__2218 (
            .O(N__16842),
            .I(N__16804));
    InMux I__2217 (
            .O(N__16841),
            .I(N__16795));
    InMux I__2216 (
            .O(N__16840),
            .I(N__16795));
    InMux I__2215 (
            .O(N__16837),
            .I(N__16795));
    InMux I__2214 (
            .O(N__16836),
            .I(N__16795));
    LocalMux I__2213 (
            .O(N__16833),
            .I(N__16792));
    InMux I__2212 (
            .O(N__16830),
            .I(N__16789));
    InMux I__2211 (
            .O(N__16827),
            .I(N__16786));
    InMux I__2210 (
            .O(N__16824),
            .I(N__16781));
    InMux I__2209 (
            .O(N__16823),
            .I(N__16781));
    CascadeMux I__2208 (
            .O(N__16822),
            .I(N__16775));
    InMux I__2207 (
            .O(N__16819),
            .I(N__16771));
    InMux I__2206 (
            .O(N__16818),
            .I(N__16768));
    Span4Mux_h I__2205 (
            .O(N__16815),
            .I(N__16765));
    Span4Mux_h I__2204 (
            .O(N__16812),
            .I(N__16756));
    LocalMux I__2203 (
            .O(N__16809),
            .I(N__16756));
    LocalMux I__2202 (
            .O(N__16804),
            .I(N__16756));
    LocalMux I__2201 (
            .O(N__16795),
            .I(N__16756));
    Span4Mux_h I__2200 (
            .O(N__16792),
            .I(N__16753));
    LocalMux I__2199 (
            .O(N__16789),
            .I(N__16746));
    LocalMux I__2198 (
            .O(N__16786),
            .I(N__16746));
    LocalMux I__2197 (
            .O(N__16781),
            .I(N__16746));
    InMux I__2196 (
            .O(N__16780),
            .I(N__16743));
    InMux I__2195 (
            .O(N__16779),
            .I(N__16738));
    InMux I__2194 (
            .O(N__16778),
            .I(N__16738));
    InMux I__2193 (
            .O(N__16775),
            .I(N__16733));
    InMux I__2192 (
            .O(N__16774),
            .I(N__16733));
    LocalMux I__2191 (
            .O(N__16771),
            .I(N__16728));
    LocalMux I__2190 (
            .O(N__16768),
            .I(N__16728));
    Span4Mux_s0_h I__2189 (
            .O(N__16765),
            .I(N__16723));
    Span4Mux_v I__2188 (
            .O(N__16756),
            .I(N__16723));
    Odrv4 I__2187 (
            .O(N__16753),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2186 (
            .O(N__16746),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2185 (
            .O(N__16743),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2184 (
            .O(N__16738),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__2183 (
            .O(N__16733),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv12 I__2182 (
            .O(N__16728),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__2181 (
            .O(N__16723),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    InMux I__2180 (
            .O(N__16708),
            .I(N__16699));
    InMux I__2179 (
            .O(N__16707),
            .I(N__16695));
    InMux I__2178 (
            .O(N__16706),
            .I(N__16692));
    InMux I__2177 (
            .O(N__16705),
            .I(N__16689));
    CascadeMux I__2176 (
            .O(N__16704),
            .I(N__16683));
    InMux I__2175 (
            .O(N__16703),
            .I(N__16675));
    InMux I__2174 (
            .O(N__16702),
            .I(N__16675));
    LocalMux I__2173 (
            .O(N__16699),
            .I(N__16672));
    InMux I__2172 (
            .O(N__16698),
            .I(N__16669));
    LocalMux I__2171 (
            .O(N__16695),
            .I(N__16666));
    LocalMux I__2170 (
            .O(N__16692),
            .I(N__16663));
    LocalMux I__2169 (
            .O(N__16689),
            .I(N__16660));
    InMux I__2168 (
            .O(N__16688),
            .I(N__16657));
    InMux I__2167 (
            .O(N__16687),
            .I(N__16654));
    InMux I__2166 (
            .O(N__16686),
            .I(N__16651));
    InMux I__2165 (
            .O(N__16683),
            .I(N__16646));
    InMux I__2164 (
            .O(N__16682),
            .I(N__16646));
    InMux I__2163 (
            .O(N__16681),
            .I(N__16643));
    InMux I__2162 (
            .O(N__16680),
            .I(N__16640));
    LocalMux I__2161 (
            .O(N__16675),
            .I(N__16633));
    Span4Mux_h I__2160 (
            .O(N__16672),
            .I(N__16633));
    LocalMux I__2159 (
            .O(N__16669),
            .I(N__16633));
    Span4Mux_v I__2158 (
            .O(N__16666),
            .I(N__16624));
    Span4Mux_v I__2157 (
            .O(N__16663),
            .I(N__16624));
    Span4Mux_v I__2156 (
            .O(N__16660),
            .I(N__16624));
    LocalMux I__2155 (
            .O(N__16657),
            .I(N__16624));
    LocalMux I__2154 (
            .O(N__16654),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__2153 (
            .O(N__16651),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__2152 (
            .O(N__16646),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__2151 (
            .O(N__16643),
            .I(this_vga_signals_M_vcounter_q_7));
    LocalMux I__2150 (
            .O(N__16640),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__2149 (
            .O(N__16633),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__2148 (
            .O(N__16624),
            .I(this_vga_signals_M_vcounter_q_7));
    InMux I__2147 (
            .O(N__16609),
            .I(N__16606));
    LocalMux I__2146 (
            .O(N__16606),
            .I(\this_vga_signals.g0_0_2 ));
    InMux I__2145 (
            .O(N__16603),
            .I(N__16598));
    InMux I__2144 (
            .O(N__16602),
            .I(N__16595));
    InMux I__2143 (
            .O(N__16601),
            .I(N__16587));
    LocalMux I__2142 (
            .O(N__16598),
            .I(N__16584));
    LocalMux I__2141 (
            .O(N__16595),
            .I(N__16581));
    InMux I__2140 (
            .O(N__16594),
            .I(N__16575));
    InMux I__2139 (
            .O(N__16593),
            .I(N__16575));
    InMux I__2138 (
            .O(N__16592),
            .I(N__16568));
    InMux I__2137 (
            .O(N__16591),
            .I(N__16568));
    InMux I__2136 (
            .O(N__16590),
            .I(N__16568));
    LocalMux I__2135 (
            .O(N__16587),
            .I(N__16558));
    Span4Mux_v I__2134 (
            .O(N__16584),
            .I(N__16558));
    Span4Mux_v I__2133 (
            .O(N__16581),
            .I(N__16558));
    InMux I__2132 (
            .O(N__16580),
            .I(N__16555));
    LocalMux I__2131 (
            .O(N__16575),
            .I(N__16550));
    LocalMux I__2130 (
            .O(N__16568),
            .I(N__16550));
    InMux I__2129 (
            .O(N__16567),
            .I(N__16547));
    InMux I__2128 (
            .O(N__16566),
            .I(N__16542));
    InMux I__2127 (
            .O(N__16565),
            .I(N__16542));
    Odrv4 I__2126 (
            .O(N__16558),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__2125 (
            .O(N__16555),
            .I(\this_vga_signals.vaddress_c2 ));
    Odrv4 I__2124 (
            .O(N__16550),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__2123 (
            .O(N__16547),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__2122 (
            .O(N__16542),
            .I(\this_vga_signals.vaddress_c2 ));
    CascadeMux I__2121 (
            .O(N__16531),
            .I(N__16528));
    InMux I__2120 (
            .O(N__16528),
            .I(N__16525));
    LocalMux I__2119 (
            .O(N__16525),
            .I(N__16522));
    Span4Mux_s2_h I__2118 (
            .O(N__16522),
            .I(N__16519));
    Odrv4 I__2117 (
            .O(N__16519),
            .I(\this_vga_signals.g0_0_3_0 ));
    SRMux I__2116 (
            .O(N__16516),
            .I(N__16511));
    SRMux I__2115 (
            .O(N__16515),
            .I(N__16508));
    SRMux I__2114 (
            .O(N__16514),
            .I(N__16505));
    LocalMux I__2113 (
            .O(N__16511),
            .I(N__16502));
    LocalMux I__2112 (
            .O(N__16508),
            .I(N__16499));
    LocalMux I__2111 (
            .O(N__16505),
            .I(N__16496));
    Span4Mux_v I__2110 (
            .O(N__16502),
            .I(N__16492));
    Span4Mux_v I__2109 (
            .O(N__16499),
            .I(N__16487));
    Span4Mux_h I__2108 (
            .O(N__16496),
            .I(N__16487));
    InMux I__2107 (
            .O(N__16495),
            .I(N__16484));
    Odrv4 I__2106 (
            .O(N__16492),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9 ));
    Odrv4 I__2105 (
            .O(N__16487),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9 ));
    LocalMux I__2104 (
            .O(N__16484),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9 ));
    CEMux I__2103 (
            .O(N__16477),
            .I(N__16474));
    LocalMux I__2102 (
            .O(N__16474),
            .I(N__16471));
    Span4Mux_h I__2101 (
            .O(N__16471),
            .I(N__16468));
    Span4Mux_h I__2100 (
            .O(N__16468),
            .I(N__16465));
    Odrv4 I__2099 (
            .O(N__16465),
            .I(\this_vga_signals.N_935_1 ));
    InMux I__2098 (
            .O(N__16462),
            .I(N__16459));
    LocalMux I__2097 (
            .O(N__16459),
            .I(N__16456));
    Span4Mux_h I__2096 (
            .O(N__16456),
            .I(N__16453));
    Odrv4 I__2095 (
            .O(N__16453),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    CascadeMux I__2094 (
            .O(N__16450),
            .I(N__16447));
    InMux I__2093 (
            .O(N__16447),
            .I(N__16444));
    LocalMux I__2092 (
            .O(N__16444),
            .I(\this_vga_signals.g0_0_0 ));
    IoInMux I__2091 (
            .O(N__16441),
            .I(N__16438));
    LocalMux I__2090 (
            .O(N__16438),
            .I(N__16435));
    Span12Mux_s9_v I__2089 (
            .O(N__16435),
            .I(N__16432));
    Odrv12 I__2088 (
            .O(N__16432),
            .I(M_vcounter_q_esr_RNIQJSA2_0_9));
    InMux I__2087 (
            .O(N__16429),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__2086 (
            .O(N__16426),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__2085 (
            .O(N__16423),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__2084 (
            .O(N__16420),
            .I(bfn_5_10_0_));
    CascadeMux I__2083 (
            .O(N__16417),
            .I(\this_vga_signals.un4_hsynclto3_0_cascade_ ));
    InMux I__2082 (
            .O(N__16414),
            .I(N__16411));
    LocalMux I__2081 (
            .O(N__16411),
            .I(this_vga_signals_un4_lvisibility_1));
    InMux I__2080 (
            .O(N__16408),
            .I(N__16404));
    CascadeMux I__2079 (
            .O(N__16407),
            .I(N__16401));
    LocalMux I__2078 (
            .O(N__16404),
            .I(N__16394));
    InMux I__2077 (
            .O(N__16401),
            .I(N__16391));
    InMux I__2076 (
            .O(N__16400),
            .I(N__16388));
    InMux I__2075 (
            .O(N__16399),
            .I(N__16382));
    InMux I__2074 (
            .O(N__16398),
            .I(N__16382));
    InMux I__2073 (
            .O(N__16397),
            .I(N__16373));
    Span4Mux_v I__2072 (
            .O(N__16394),
            .I(N__16368));
    LocalMux I__2071 (
            .O(N__16391),
            .I(N__16368));
    LocalMux I__2070 (
            .O(N__16388),
            .I(N__16365));
    InMux I__2069 (
            .O(N__16387),
            .I(N__16362));
    LocalMux I__2068 (
            .O(N__16382),
            .I(N__16359));
    InMux I__2067 (
            .O(N__16381),
            .I(N__16356));
    InMux I__2066 (
            .O(N__16380),
            .I(N__16351));
    InMux I__2065 (
            .O(N__16379),
            .I(N__16351));
    InMux I__2064 (
            .O(N__16378),
            .I(N__16346));
    InMux I__2063 (
            .O(N__16377),
            .I(N__16346));
    InMux I__2062 (
            .O(N__16376),
            .I(N__16343));
    LocalMux I__2061 (
            .O(N__16373),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__2060 (
            .O(N__16368),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__2059 (
            .O(N__16365),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__2058 (
            .O(N__16362),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__2057 (
            .O(N__16359),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__2056 (
            .O(N__16356),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__2055 (
            .O(N__16351),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__2054 (
            .O(N__16346),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__2053 (
            .O(N__16343),
            .I(this_vga_signals_M_vcounter_q_8));
    InMux I__2052 (
            .O(N__16324),
            .I(N__16321));
    LocalMux I__2051 (
            .O(N__16321),
            .I(N__16317));
    InMux I__2050 (
            .O(N__16320),
            .I(N__16314));
    Span4Mux_h I__2049 (
            .O(N__16317),
            .I(N__16308));
    LocalMux I__2048 (
            .O(N__16314),
            .I(N__16308));
    InMux I__2047 (
            .O(N__16313),
            .I(N__16305));
    Odrv4 I__2046 (
            .O(N__16308),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    LocalMux I__2045 (
            .O(N__16305),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    CEMux I__2044 (
            .O(N__16300),
            .I(N__16273));
    CEMux I__2043 (
            .O(N__16299),
            .I(N__16273));
    CEMux I__2042 (
            .O(N__16298),
            .I(N__16273));
    CEMux I__2041 (
            .O(N__16297),
            .I(N__16273));
    CEMux I__2040 (
            .O(N__16296),
            .I(N__16273));
    CEMux I__2039 (
            .O(N__16295),
            .I(N__16273));
    CEMux I__2038 (
            .O(N__16294),
            .I(N__16273));
    CEMux I__2037 (
            .O(N__16293),
            .I(N__16273));
    CEMux I__2036 (
            .O(N__16292),
            .I(N__16273));
    GlobalMux I__2035 (
            .O(N__16273),
            .I(N__16270));
    gio2CtrlBuf I__2034 (
            .O(N__16270),
            .I(\this_vga_signals.N_935_0_g ));
    InMux I__2033 (
            .O(N__16267),
            .I(N__16264));
    LocalMux I__2032 (
            .O(N__16264),
            .I(N__16251));
    SRMux I__2031 (
            .O(N__16263),
            .I(N__16228));
    SRMux I__2030 (
            .O(N__16262),
            .I(N__16228));
    SRMux I__2029 (
            .O(N__16261),
            .I(N__16228));
    SRMux I__2028 (
            .O(N__16260),
            .I(N__16228));
    SRMux I__2027 (
            .O(N__16259),
            .I(N__16228));
    SRMux I__2026 (
            .O(N__16258),
            .I(N__16228));
    SRMux I__2025 (
            .O(N__16257),
            .I(N__16228));
    SRMux I__2024 (
            .O(N__16256),
            .I(N__16228));
    SRMux I__2023 (
            .O(N__16255),
            .I(N__16228));
    SRMux I__2022 (
            .O(N__16254),
            .I(N__16228));
    Glb2LocalMux I__2021 (
            .O(N__16251),
            .I(N__16228));
    GlobalMux I__2020 (
            .O(N__16228),
            .I(N__16225));
    gio2CtrlBuf I__2019 (
            .O(N__16225),
            .I(\this_vga_signals.N_1212_g ));
    InMux I__2018 (
            .O(N__16222),
            .I(N__16219));
    LocalMux I__2017 (
            .O(N__16219),
            .I(N__16216));
    Odrv4 I__2016 (
            .O(N__16216),
            .I(\this_vga_signals.un4_hsynclto7_0 ));
    InMux I__2015 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__2014 (
            .O(N__16210),
            .I(N__16207));
    Span4Mux_v I__2013 (
            .O(N__16207),
            .I(N__16204));
    Odrv4 I__2012 (
            .O(N__16204),
            .I(\this_vga_signals.un4_hsynclt9 ));
    CascadeMux I__2011 (
            .O(N__16201),
            .I(\this_vga_signals.if_N_8_i_0_cascade_ ));
    CascadeMux I__2010 (
            .O(N__16198),
            .I(\this_vga_signals.if_N_9_0_0_cascade_ ));
    InMux I__2009 (
            .O(N__16195),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__2008 (
            .O(N__16192),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__2007 (
            .O(N__16189),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__2006 (
            .O(N__16186),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    CascadeMux I__2005 (
            .O(N__16183),
            .I(\this_vga_signals.r_N_4_mux_cascade_ ));
    InMux I__2004 (
            .O(N__16180),
            .I(N__16176));
    InMux I__2003 (
            .O(N__16179),
            .I(N__16173));
    LocalMux I__2002 (
            .O(N__16176),
            .I(\this_vga_signals.N_24_0 ));
    LocalMux I__2001 (
            .O(N__16173),
            .I(\this_vga_signals.N_24_0 ));
    InMux I__2000 (
            .O(N__16168),
            .I(N__16165));
    LocalMux I__1999 (
            .O(N__16165),
            .I(\this_vga_signals.r_N_4_mux ));
    InMux I__1998 (
            .O(N__16162),
            .I(N__16157));
    InMux I__1997 (
            .O(N__16161),
            .I(N__16151));
    InMux I__1996 (
            .O(N__16160),
            .I(N__16148));
    LocalMux I__1995 (
            .O(N__16157),
            .I(N__16145));
    InMux I__1994 (
            .O(N__16156),
            .I(N__16140));
    InMux I__1993 (
            .O(N__16155),
            .I(N__16140));
    InMux I__1992 (
            .O(N__16154),
            .I(N__16137));
    LocalMux I__1991 (
            .O(N__16151),
            .I(N__16134));
    LocalMux I__1990 (
            .O(N__16148),
            .I(N__16130));
    Span4Mux_v I__1989 (
            .O(N__16145),
            .I(N__16123));
    LocalMux I__1988 (
            .O(N__16140),
            .I(N__16123));
    LocalMux I__1987 (
            .O(N__16137),
            .I(N__16123));
    Span4Mux_v I__1986 (
            .O(N__16134),
            .I(N__16120));
    InMux I__1985 (
            .O(N__16133),
            .I(N__16117));
    Span4Mux_v I__1984 (
            .O(N__16130),
            .I(N__16114));
    Span4Mux_h I__1983 (
            .O(N__16123),
            .I(N__16111));
    Odrv4 I__1982 (
            .O(N__16120),
            .I(\this_vga_signals.N_32_0 ));
    LocalMux I__1981 (
            .O(N__16117),
            .I(\this_vga_signals.N_32_0 ));
    Odrv4 I__1980 (
            .O(N__16114),
            .I(\this_vga_signals.N_32_0 ));
    Odrv4 I__1979 (
            .O(N__16111),
            .I(\this_vga_signals.N_32_0 ));
    CascadeMux I__1978 (
            .O(N__16102),
            .I(\this_vga_signals.N_24_0_2_cascade_ ));
    InMux I__1977 (
            .O(N__16099),
            .I(N__16093));
    InMux I__1976 (
            .O(N__16098),
            .I(N__16090));
    InMux I__1975 (
            .O(N__16097),
            .I(N__16087));
    InMux I__1974 (
            .O(N__16096),
            .I(N__16084));
    LocalMux I__1973 (
            .O(N__16093),
            .I(\this_vga_signals.mult1_un40_sum_c2_0 ));
    LocalMux I__1972 (
            .O(N__16090),
            .I(\this_vga_signals.mult1_un40_sum_c2_0 ));
    LocalMux I__1971 (
            .O(N__16087),
            .I(\this_vga_signals.mult1_un40_sum_c2_0 ));
    LocalMux I__1970 (
            .O(N__16084),
            .I(\this_vga_signals.mult1_un40_sum_c2_0 ));
    InMux I__1969 (
            .O(N__16075),
            .I(N__16072));
    LocalMux I__1968 (
            .O(N__16072),
            .I(N__16068));
    InMux I__1967 (
            .O(N__16071),
            .I(N__16065));
    Odrv4 I__1966 (
            .O(N__16068),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1 ));
    LocalMux I__1965 (
            .O(N__16065),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1 ));
    InMux I__1964 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__1963 (
            .O(N__16057),
            .I(N__16052));
    InMux I__1962 (
            .O(N__16056),
            .I(N__16047));
    InMux I__1961 (
            .O(N__16055),
            .I(N__16047));
    Span4Mux_v I__1960 (
            .O(N__16052),
            .I(N__16041));
    LocalMux I__1959 (
            .O(N__16047),
            .I(N__16041));
    InMux I__1958 (
            .O(N__16046),
            .I(N__16038));
    Span4Mux_h I__1957 (
            .O(N__16041),
            .I(N__16035));
    LocalMux I__1956 (
            .O(N__16038),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_0 ));
    Odrv4 I__1955 (
            .O(N__16035),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_0 ));
    CascadeMux I__1954 (
            .O(N__16030),
            .I(\this_vga_signals.g0_23_cascade_ ));
    InMux I__1953 (
            .O(N__16027),
            .I(N__16020));
    InMux I__1952 (
            .O(N__16026),
            .I(N__16015));
    InMux I__1951 (
            .O(N__16025),
            .I(N__16015));
    InMux I__1950 (
            .O(N__16024),
            .I(N__16010));
    InMux I__1949 (
            .O(N__16023),
            .I(N__16010));
    LocalMux I__1948 (
            .O(N__16020),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ));
    LocalMux I__1947 (
            .O(N__16015),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ));
    LocalMux I__1946 (
            .O(N__16010),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ));
    CascadeMux I__1945 (
            .O(N__16003),
            .I(N__16000));
    InMux I__1944 (
            .O(N__16000),
            .I(N__15997));
    LocalMux I__1943 (
            .O(N__15997),
            .I(\this_vga_signals.g0_1_0_0 ));
    InMux I__1942 (
            .O(N__15994),
            .I(N__15991));
    LocalMux I__1941 (
            .O(N__15991),
            .I(\this_vga_signals.g1_0_0 ));
    InMux I__1940 (
            .O(N__15988),
            .I(N__15985));
    LocalMux I__1939 (
            .O(N__15985),
            .I(\this_vga_signals.g0_0_2_0 ));
    InMux I__1938 (
            .O(N__15982),
            .I(N__15979));
    LocalMux I__1937 (
            .O(N__15979),
            .I(N__15976));
    Odrv12 I__1936 (
            .O(N__15976),
            .I(\this_vga_signals.un2_hsynclt7 ));
    IoInMux I__1935 (
            .O(N__15973),
            .I(N__15970));
    LocalMux I__1934 (
            .O(N__15970),
            .I(N__15967));
    IoSpan4Mux I__1933 (
            .O(N__15967),
            .I(N__15964));
    Sp12to4 I__1932 (
            .O(N__15964),
            .I(N__15961));
    Span12Mux_s6_v I__1931 (
            .O(N__15961),
            .I(N__15958));
    Odrv12 I__1930 (
            .O(N__15958),
            .I(this_vga_signals_hsync_1_i));
    IoInMux I__1929 (
            .O(N__15955),
            .I(N__15952));
    LocalMux I__1928 (
            .O(N__15952),
            .I(N__15949));
    Span4Mux_s3_h I__1927 (
            .O(N__15949),
            .I(N__15946));
    Span4Mux_v I__1926 (
            .O(N__15946),
            .I(N__15943));
    Span4Mux_v I__1925 (
            .O(N__15943),
            .I(N__15940));
    Odrv4 I__1924 (
            .O(N__15940),
            .I(rgb_c_5));
    CascadeMux I__1923 (
            .O(N__15937),
            .I(\this_vga_signals.r_N_4_mux_1_cascade_ ));
    InMux I__1922 (
            .O(N__15934),
            .I(N__15931));
    LocalMux I__1921 (
            .O(N__15931),
            .I(N__15928));
    Odrv4 I__1920 (
            .O(N__15928),
            .I(\this_vga_signals.N_24_0_1 ));
    CascadeMux I__1919 (
            .O(N__15925),
            .I(\this_vga_signals.un2_hsynclt6_0_cascade_ ));
    InMux I__1918 (
            .O(N__15922),
            .I(N__15919));
    LocalMux I__1917 (
            .O(N__15919),
            .I(N__15914));
    InMux I__1916 (
            .O(N__15918),
            .I(N__15911));
    InMux I__1915 (
            .O(N__15917),
            .I(N__15908));
    Odrv4 I__1914 (
            .O(N__15914),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    LocalMux I__1913 (
            .O(N__15911),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    LocalMux I__1912 (
            .O(N__15908),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    InMux I__1911 (
            .O(N__15901),
            .I(N__15898));
    LocalMux I__1910 (
            .O(N__15898),
            .I(N__15895));
    Odrv4 I__1909 (
            .O(N__15895),
            .I(\this_vga_signals.r_N_4_mux_0 ));
    CascadeMux I__1908 (
            .O(N__15892),
            .I(\this_vga_signals.N_24_0_0_cascade_ ));
    InMux I__1907 (
            .O(N__15889),
            .I(N__15883));
    InMux I__1906 (
            .O(N__15888),
            .I(N__15883));
    LocalMux I__1905 (
            .O(N__15883),
            .I(\this_vga_signals.N_4_2_0 ));
    InMux I__1904 (
            .O(N__15880),
            .I(N__15877));
    LocalMux I__1903 (
            .O(N__15877),
            .I(N__15873));
    InMux I__1902 (
            .O(N__15876),
            .I(N__15870));
    Span4Mux_v I__1901 (
            .O(N__15873),
            .I(N__15864));
    LocalMux I__1900 (
            .O(N__15870),
            .I(N__15864));
    InMux I__1899 (
            .O(N__15869),
            .I(N__15861));
    Odrv4 I__1898 (
            .O(N__15864),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    LocalMux I__1897 (
            .O(N__15861),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    InMux I__1896 (
            .O(N__15856),
            .I(N__15853));
    LocalMux I__1895 (
            .O(N__15853),
            .I(N__15850));
    Span4Mux_s3_h I__1894 (
            .O(N__15850),
            .I(N__15847));
    Odrv4 I__1893 (
            .O(N__15847),
            .I(\this_vga_signals.g0_0_i_a5_1_0 ));
    InMux I__1892 (
            .O(N__15844),
            .I(N__15841));
    LocalMux I__1891 (
            .O(N__15841),
            .I(N__15834));
    InMux I__1890 (
            .O(N__15840),
            .I(N__15831));
    CascadeMux I__1889 (
            .O(N__15839),
            .I(N__15828));
    InMux I__1888 (
            .O(N__15838),
            .I(N__15825));
    InMux I__1887 (
            .O(N__15837),
            .I(N__15818));
    Span4Mux_h I__1886 (
            .O(N__15834),
            .I(N__15815));
    LocalMux I__1885 (
            .O(N__15831),
            .I(N__15812));
    InMux I__1884 (
            .O(N__15828),
            .I(N__15809));
    LocalMux I__1883 (
            .O(N__15825),
            .I(N__15806));
    InMux I__1882 (
            .O(N__15824),
            .I(N__15797));
    InMux I__1881 (
            .O(N__15823),
            .I(N__15797));
    InMux I__1880 (
            .O(N__15822),
            .I(N__15797));
    InMux I__1879 (
            .O(N__15821),
            .I(N__15797));
    LocalMux I__1878 (
            .O(N__15818),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__1877 (
            .O(N__15815),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv12 I__1876 (
            .O(N__15812),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1875 (
            .O(N__15809),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    Odrv4 I__1874 (
            .O(N__15806),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__1873 (
            .O(N__15797),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    InMux I__1872 (
            .O(N__15784),
            .I(N__15779));
    InMux I__1871 (
            .O(N__15783),
            .I(N__15774));
    InMux I__1870 (
            .O(N__15782),
            .I(N__15774));
    LocalMux I__1869 (
            .O(N__15779),
            .I(N__15769));
    LocalMux I__1868 (
            .O(N__15774),
            .I(N__15766));
    CascadeMux I__1867 (
            .O(N__15773),
            .I(N__15758));
    InMux I__1866 (
            .O(N__15772),
            .I(N__15754));
    Span4Mux_h I__1865 (
            .O(N__15769),
            .I(N__15751));
    Span4Mux_h I__1864 (
            .O(N__15766),
            .I(N__15748));
    InMux I__1863 (
            .O(N__15765),
            .I(N__15745));
    InMux I__1862 (
            .O(N__15764),
            .I(N__15732));
    InMux I__1861 (
            .O(N__15763),
            .I(N__15732));
    InMux I__1860 (
            .O(N__15762),
            .I(N__15732));
    InMux I__1859 (
            .O(N__15761),
            .I(N__15732));
    InMux I__1858 (
            .O(N__15758),
            .I(N__15732));
    InMux I__1857 (
            .O(N__15757),
            .I(N__15732));
    LocalMux I__1856 (
            .O(N__15754),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__1855 (
            .O(N__15751),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    Odrv4 I__1854 (
            .O(N__15748),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__1853 (
            .O(N__15745),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__1852 (
            .O(N__15732),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    InMux I__1851 (
            .O(N__15721),
            .I(N__15718));
    LocalMux I__1850 (
            .O(N__15718),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    CascadeMux I__1849 (
            .O(N__15715),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ));
    InMux I__1848 (
            .O(N__15712),
            .I(N__15709));
    LocalMux I__1847 (
            .O(N__15709),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_0_0 ));
    CascadeMux I__1846 (
            .O(N__15706),
            .I(\this_vga_signals.vvisibility_i_o2_1_cascade_ ));
    InMux I__1845 (
            .O(N__15703),
            .I(N__15700));
    LocalMux I__1844 (
            .O(N__15700),
            .I(N__15696));
    InMux I__1843 (
            .O(N__15699),
            .I(N__15693));
    Odrv4 I__1842 (
            .O(N__15696),
            .I(\this_vga_signals.vaddress_m2_e_1 ));
    LocalMux I__1841 (
            .O(N__15693),
            .I(\this_vga_signals.vaddress_m2_e_1 ));
    InMux I__1840 (
            .O(N__15688),
            .I(N__15684));
    InMux I__1839 (
            .O(N__15687),
            .I(N__15681));
    LocalMux I__1838 (
            .O(N__15684),
            .I(N__15674));
    LocalMux I__1837 (
            .O(N__15681),
            .I(N__15674));
    InMux I__1836 (
            .O(N__15680),
            .I(N__15667));
    InMux I__1835 (
            .O(N__15679),
            .I(N__15667));
    Span4Mux_v I__1834 (
            .O(N__15674),
            .I(N__15664));
    InMux I__1833 (
            .O(N__15673),
            .I(N__15661));
    InMux I__1832 (
            .O(N__15672),
            .I(N__15657));
    LocalMux I__1831 (
            .O(N__15667),
            .I(N__15654));
    Span4Mux_v I__1830 (
            .O(N__15664),
            .I(N__15649));
    LocalMux I__1829 (
            .O(N__15661),
            .I(N__15649));
    InMux I__1828 (
            .O(N__15660),
            .I(N__15646));
    LocalMux I__1827 (
            .O(N__15657),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv12 I__1826 (
            .O(N__15654),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv4 I__1825 (
            .O(N__15649),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__1824 (
            .O(N__15646),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    InMux I__1823 (
            .O(N__15637),
            .I(N__15634));
    LocalMux I__1822 (
            .O(N__15634),
            .I(N__15628));
    InMux I__1821 (
            .O(N__15633),
            .I(N__15622));
    InMux I__1820 (
            .O(N__15632),
            .I(N__15622));
    InMux I__1819 (
            .O(N__15631),
            .I(N__15617));
    Span4Mux_v I__1818 (
            .O(N__15628),
            .I(N__15614));
    InMux I__1817 (
            .O(N__15627),
            .I(N__15611));
    LocalMux I__1816 (
            .O(N__15622),
            .I(N__15606));
    InMux I__1815 (
            .O(N__15621),
            .I(N__15603));
    InMux I__1814 (
            .O(N__15620),
            .I(N__15600));
    LocalMux I__1813 (
            .O(N__15617),
            .I(N__15594));
    IoSpan4Mux I__1812 (
            .O(N__15614),
            .I(N__15591));
    LocalMux I__1811 (
            .O(N__15611),
            .I(N__15588));
    InMux I__1810 (
            .O(N__15610),
            .I(N__15583));
    InMux I__1809 (
            .O(N__15609),
            .I(N__15583));
    Span4Mux_s2_h I__1808 (
            .O(N__15606),
            .I(N__15580));
    LocalMux I__1807 (
            .O(N__15603),
            .I(N__15577));
    LocalMux I__1806 (
            .O(N__15600),
            .I(N__15573));
    InMux I__1805 (
            .O(N__15599),
            .I(N__15570));
    InMux I__1804 (
            .O(N__15598),
            .I(N__15565));
    InMux I__1803 (
            .O(N__15597),
            .I(N__15565));
    Span4Mux_v I__1802 (
            .O(N__15594),
            .I(N__15558));
    Span4Mux_s2_h I__1801 (
            .O(N__15591),
            .I(N__15558));
    Span4Mux_s2_h I__1800 (
            .O(N__15588),
            .I(N__15558));
    LocalMux I__1799 (
            .O(N__15583),
            .I(N__15551));
    Span4Mux_h I__1798 (
            .O(N__15580),
            .I(N__15551));
    Span4Mux_s2_h I__1797 (
            .O(N__15577),
            .I(N__15551));
    InMux I__1796 (
            .O(N__15576),
            .I(N__15547));
    Span4Mux_s2_h I__1795 (
            .O(N__15573),
            .I(N__15544));
    LocalMux I__1794 (
            .O(N__15570),
            .I(N__15541));
    LocalMux I__1793 (
            .O(N__15565),
            .I(N__15534));
    Sp12to4 I__1792 (
            .O(N__15558),
            .I(N__15534));
    Sp12to4 I__1791 (
            .O(N__15551),
            .I(N__15534));
    InMux I__1790 (
            .O(N__15550),
            .I(N__15531));
    LocalMux I__1789 (
            .O(N__15547),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1788 (
            .O(N__15544),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__1787 (
            .O(N__15541),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv12 I__1786 (
            .O(N__15534),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__1785 (
            .O(N__15531),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    CascadeMux I__1784 (
            .O(N__15520),
            .I(N__15509));
    CascadeMux I__1783 (
            .O(N__15519),
            .I(N__15506));
    CascadeMux I__1782 (
            .O(N__15518),
            .I(N__15502));
    CascadeMux I__1781 (
            .O(N__15517),
            .I(N__15499));
    CascadeMux I__1780 (
            .O(N__15516),
            .I(N__15495));
    CascadeMux I__1779 (
            .O(N__15515),
            .I(N__15492));
    CascadeMux I__1778 (
            .O(N__15514),
            .I(N__15487));
    CascadeMux I__1777 (
            .O(N__15513),
            .I(N__15484));
    CascadeMux I__1776 (
            .O(N__15512),
            .I(N__15481));
    InMux I__1775 (
            .O(N__15509),
            .I(N__15477));
    InMux I__1774 (
            .O(N__15506),
            .I(N__15473));
    InMux I__1773 (
            .O(N__15505),
            .I(N__15470));
    InMux I__1772 (
            .O(N__15502),
            .I(N__15467));
    InMux I__1771 (
            .O(N__15499),
            .I(N__15458));
    InMux I__1770 (
            .O(N__15498),
            .I(N__15458));
    InMux I__1769 (
            .O(N__15495),
            .I(N__15458));
    InMux I__1768 (
            .O(N__15492),
            .I(N__15458));
    InMux I__1767 (
            .O(N__15491),
            .I(N__15455));
    InMux I__1766 (
            .O(N__15490),
            .I(N__15452));
    InMux I__1765 (
            .O(N__15487),
            .I(N__15449));
    InMux I__1764 (
            .O(N__15484),
            .I(N__15444));
    InMux I__1763 (
            .O(N__15481),
            .I(N__15444));
    InMux I__1762 (
            .O(N__15480),
            .I(N__15441));
    LocalMux I__1761 (
            .O(N__15477),
            .I(N__15438));
    InMux I__1760 (
            .O(N__15476),
            .I(N__15435));
    LocalMux I__1759 (
            .O(N__15473),
            .I(N__15430));
    LocalMux I__1758 (
            .O(N__15470),
            .I(N__15430));
    LocalMux I__1757 (
            .O(N__15467),
            .I(N__15425));
    LocalMux I__1756 (
            .O(N__15458),
            .I(N__15425));
    LocalMux I__1755 (
            .O(N__15455),
            .I(N__15417));
    LocalMux I__1754 (
            .O(N__15452),
            .I(N__15417));
    LocalMux I__1753 (
            .O(N__15449),
            .I(N__15412));
    LocalMux I__1752 (
            .O(N__15444),
            .I(N__15412));
    LocalMux I__1751 (
            .O(N__15441),
            .I(N__15401));
    Span4Mux_s1_h I__1750 (
            .O(N__15438),
            .I(N__15401));
    LocalMux I__1749 (
            .O(N__15435),
            .I(N__15401));
    Span4Mux_v I__1748 (
            .O(N__15430),
            .I(N__15401));
    Span4Mux_v I__1747 (
            .O(N__15425),
            .I(N__15401));
    InMux I__1746 (
            .O(N__15424),
            .I(N__15396));
    InMux I__1745 (
            .O(N__15423),
            .I(N__15393));
    InMux I__1744 (
            .O(N__15422),
            .I(N__15390));
    Span4Mux_v I__1743 (
            .O(N__15417),
            .I(N__15387));
    Span4Mux_v I__1742 (
            .O(N__15412),
            .I(N__15384));
    Span4Mux_v I__1741 (
            .O(N__15401),
            .I(N__15381));
    InMux I__1740 (
            .O(N__15400),
            .I(N__15377));
    CascadeMux I__1739 (
            .O(N__15399),
            .I(N__15374));
    LocalMux I__1738 (
            .O(N__15396),
            .I(N__15369));
    LocalMux I__1737 (
            .O(N__15393),
            .I(N__15369));
    LocalMux I__1736 (
            .O(N__15390),
            .I(N__15360));
    Span4Mux_s1_h I__1735 (
            .O(N__15387),
            .I(N__15360));
    Span4Mux_v I__1734 (
            .O(N__15384),
            .I(N__15360));
    Span4Mux_s1_h I__1733 (
            .O(N__15381),
            .I(N__15360));
    InMux I__1732 (
            .O(N__15380),
            .I(N__15357));
    LocalMux I__1731 (
            .O(N__15377),
            .I(N__15354));
    InMux I__1730 (
            .O(N__15374),
            .I(N__15351));
    Odrv12 I__1729 (
            .O(N__15369),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__1728 (
            .O(N__15360),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1727 (
            .O(N__15357),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__1726 (
            .O(N__15354),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__1725 (
            .O(N__15351),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    InMux I__1724 (
            .O(N__15340),
            .I(N__15336));
    InMux I__1723 (
            .O(N__15339),
            .I(N__15332));
    LocalMux I__1722 (
            .O(N__15336),
            .I(N__15329));
    InMux I__1721 (
            .O(N__15335),
            .I(N__15326));
    LocalMux I__1720 (
            .O(N__15332),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    Odrv12 I__1719 (
            .O(N__15329),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__1718 (
            .O(N__15326),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__1717 (
            .O(N__15319),
            .I(\this_vga_signals.N_822_0_cascade_ ));
    InMux I__1716 (
            .O(N__15316),
            .I(N__15308));
    InMux I__1715 (
            .O(N__15315),
            .I(N__15308));
    CascadeMux I__1714 (
            .O(N__15314),
            .I(N__15302));
    CascadeMux I__1713 (
            .O(N__15313),
            .I(N__15299));
    LocalMux I__1712 (
            .O(N__15308),
            .I(N__15296));
    InMux I__1711 (
            .O(N__15307),
            .I(N__15293));
    InMux I__1710 (
            .O(N__15306),
            .I(N__15290));
    InMux I__1709 (
            .O(N__15305),
            .I(N__15285));
    InMux I__1708 (
            .O(N__15302),
            .I(N__15285));
    InMux I__1707 (
            .O(N__15299),
            .I(N__15282));
    Odrv4 I__1706 (
            .O(N__15296),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1705 (
            .O(N__15293),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1704 (
            .O(N__15290),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1703 (
            .O(N__15285),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    LocalMux I__1702 (
            .O(N__15282),
            .I(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ));
    InMux I__1701 (
            .O(N__15271),
            .I(N__15265));
    CascadeMux I__1700 (
            .O(N__15270),
            .I(N__15257));
    InMux I__1699 (
            .O(N__15269),
            .I(N__15248));
    InMux I__1698 (
            .O(N__15268),
            .I(N__15248));
    LocalMux I__1697 (
            .O(N__15265),
            .I(N__15245));
    InMux I__1696 (
            .O(N__15264),
            .I(N__15242));
    InMux I__1695 (
            .O(N__15263),
            .I(N__15235));
    InMux I__1694 (
            .O(N__15262),
            .I(N__15235));
    InMux I__1693 (
            .O(N__15261),
            .I(N__15235));
    InMux I__1692 (
            .O(N__15260),
            .I(N__15232));
    InMux I__1691 (
            .O(N__15257),
            .I(N__15225));
    InMux I__1690 (
            .O(N__15256),
            .I(N__15225));
    InMux I__1689 (
            .O(N__15255),
            .I(N__15225));
    InMux I__1688 (
            .O(N__15254),
            .I(N__15220));
    InMux I__1687 (
            .O(N__15253),
            .I(N__15220));
    LocalMux I__1686 (
            .O(N__15248),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__1685 (
            .O(N__15245),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1684 (
            .O(N__15242),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1683 (
            .O(N__15235),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1682 (
            .O(N__15232),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1681 (
            .O(N__15225),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__1680 (
            .O(N__15220),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    InMux I__1679 (
            .O(N__15205),
            .I(N__15202));
    LocalMux I__1678 (
            .O(N__15202),
            .I(N__15195));
    InMux I__1677 (
            .O(N__15201),
            .I(N__15192));
    CascadeMux I__1676 (
            .O(N__15200),
            .I(N__15189));
    CascadeMux I__1675 (
            .O(N__15199),
            .I(N__15186));
    InMux I__1674 (
            .O(N__15198),
            .I(N__15180));
    Span4Mux_s3_h I__1673 (
            .O(N__15195),
            .I(N__15177));
    LocalMux I__1672 (
            .O(N__15192),
            .I(N__15174));
    InMux I__1671 (
            .O(N__15189),
            .I(N__15171));
    InMux I__1670 (
            .O(N__15186),
            .I(N__15168));
    InMux I__1669 (
            .O(N__15185),
            .I(N__15165));
    InMux I__1668 (
            .O(N__15184),
            .I(N__15162));
    InMux I__1667 (
            .O(N__15183),
            .I(N__15159));
    LocalMux I__1666 (
            .O(N__15180),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    Odrv4 I__1665 (
            .O(N__15177),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    Odrv4 I__1664 (
            .O(N__15174),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1663 (
            .O(N__15171),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1662 (
            .O(N__15168),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1661 (
            .O(N__15165),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1660 (
            .O(N__15162),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    LocalMux I__1659 (
            .O(N__15159),
            .I(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ));
    InMux I__1658 (
            .O(N__15142),
            .I(N__15133));
    InMux I__1657 (
            .O(N__15141),
            .I(N__15128));
    InMux I__1656 (
            .O(N__15140),
            .I(N__15128));
    InMux I__1655 (
            .O(N__15139),
            .I(N__15125));
    InMux I__1654 (
            .O(N__15138),
            .I(N__15118));
    InMux I__1653 (
            .O(N__15137),
            .I(N__15118));
    InMux I__1652 (
            .O(N__15136),
            .I(N__15118));
    LocalMux I__1651 (
            .O(N__15133),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1650 (
            .O(N__15128),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1649 (
            .O(N__15125),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    LocalMux I__1648 (
            .O(N__15118),
            .I(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ));
    CascadeMux I__1647 (
            .O(N__15109),
            .I(N__15106));
    InMux I__1646 (
            .O(N__15106),
            .I(N__15103));
    LocalMux I__1645 (
            .O(N__15103),
            .I(N__15100));
    Span4Mux_s3_h I__1644 (
            .O(N__15100),
            .I(N__15097));
    Odrv4 I__1643 (
            .O(N__15097),
            .I(\this_vga_signals.mult1_un40_sum_ac0_0_0 ));
    IoInMux I__1642 (
            .O(N__15094),
            .I(N__15091));
    LocalMux I__1641 (
            .O(N__15091),
            .I(N__15088));
    Span4Mux_s2_h I__1640 (
            .O(N__15088),
            .I(N__15085));
    Odrv4 I__1639 (
            .O(N__15085),
            .I(rgb_c_2));
    InMux I__1638 (
            .O(N__15082),
            .I(N__15079));
    LocalMux I__1637 (
            .O(N__15079),
            .I(N__15076));
    Odrv4 I__1636 (
            .O(N__15076),
            .I(\this_vga_signals.vsync_1_0_a2_3 ));
    CascadeMux I__1635 (
            .O(N__15073),
            .I(N__15070));
    InMux I__1634 (
            .O(N__15070),
            .I(N__15067));
    LocalMux I__1633 (
            .O(N__15067),
            .I(\this_vga_signals.vsync_1_0_a2_4 ));
    IoInMux I__1632 (
            .O(N__15064),
            .I(N__15061));
    LocalMux I__1631 (
            .O(N__15061),
            .I(N__15058));
    Span12Mux_s11_v I__1630 (
            .O(N__15058),
            .I(N__15055));
    Odrv12 I__1629 (
            .O(N__15055),
            .I(this_vga_signals_vsync_1_i));
    InMux I__1628 (
            .O(N__15052),
            .I(N__15049));
    LocalMux I__1627 (
            .O(N__15049),
            .I(N__15046));
    Odrv4 I__1626 (
            .O(N__15046),
            .I(\this_vga_signals.if_N_6_0 ));
    CascadeMux I__1625 (
            .O(N__15043),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ));
    CascadeMux I__1624 (
            .O(N__15040),
            .I(N__15037));
    InMux I__1623 (
            .O(N__15037),
            .I(N__15034));
    LocalMux I__1622 (
            .O(N__15034),
            .I(\this_vga_signals.mult1_un75_sum_axb2_0 ));
    IoInMux I__1621 (
            .O(N__15031),
            .I(N__15028));
    LocalMux I__1620 (
            .O(N__15028),
            .I(N__15025));
    Span4Mux_s2_h I__1619 (
            .O(N__15025),
            .I(N__15022));
    Span4Mux_v I__1618 (
            .O(N__15022),
            .I(N__15019));
    Span4Mux_v I__1617 (
            .O(N__15019),
            .I(N__15016));
    Odrv4 I__1616 (
            .O(N__15016),
            .I(rgb_c_3));
    InMux I__1615 (
            .O(N__15013),
            .I(N__15009));
    InMux I__1614 (
            .O(N__15012),
            .I(N__15003));
    LocalMux I__1613 (
            .O(N__15009),
            .I(N__15000));
    InMux I__1612 (
            .O(N__15008),
            .I(N__14995));
    InMux I__1611 (
            .O(N__15007),
            .I(N__14995));
    InMux I__1610 (
            .O(N__15006),
            .I(N__14992));
    LocalMux I__1609 (
            .O(N__15003),
            .I(N__14989));
    Odrv4 I__1608 (
            .O(N__15000),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1 ));
    LocalMux I__1607 (
            .O(N__14995),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1 ));
    LocalMux I__1606 (
            .O(N__14992),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1 ));
    Odrv4 I__1605 (
            .O(N__14989),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1_1 ));
    CascadeMux I__1604 (
            .O(N__14980),
            .I(N__14975));
    InMux I__1603 (
            .O(N__14979),
            .I(N__14970));
    InMux I__1602 (
            .O(N__14978),
            .I(N__14966));
    InMux I__1601 (
            .O(N__14975),
            .I(N__14963));
    InMux I__1600 (
            .O(N__14974),
            .I(N__14955));
    CascadeMux I__1599 (
            .O(N__14973),
            .I(N__14947));
    LocalMux I__1598 (
            .O(N__14970),
            .I(N__14944));
    InMux I__1597 (
            .O(N__14969),
            .I(N__14941));
    LocalMux I__1596 (
            .O(N__14966),
            .I(N__14938));
    LocalMux I__1595 (
            .O(N__14963),
            .I(N__14935));
    InMux I__1594 (
            .O(N__14962),
            .I(N__14930));
    InMux I__1593 (
            .O(N__14961),
            .I(N__14930));
    InMux I__1592 (
            .O(N__14960),
            .I(N__14927));
    InMux I__1591 (
            .O(N__14959),
            .I(N__14922));
    InMux I__1590 (
            .O(N__14958),
            .I(N__14922));
    LocalMux I__1589 (
            .O(N__14955),
            .I(N__14919));
    InMux I__1588 (
            .O(N__14954),
            .I(N__14916));
    InMux I__1587 (
            .O(N__14953),
            .I(N__14911));
    InMux I__1586 (
            .O(N__14952),
            .I(N__14911));
    InMux I__1585 (
            .O(N__14951),
            .I(N__14904));
    InMux I__1584 (
            .O(N__14950),
            .I(N__14904));
    InMux I__1583 (
            .O(N__14947),
            .I(N__14904));
    Span4Mux_v I__1582 (
            .O(N__14944),
            .I(N__14891));
    LocalMux I__1581 (
            .O(N__14941),
            .I(N__14891));
    Span4Mux_h I__1580 (
            .O(N__14938),
            .I(N__14891));
    Span4Mux_v I__1579 (
            .O(N__14935),
            .I(N__14891));
    LocalMux I__1578 (
            .O(N__14930),
            .I(N__14891));
    LocalMux I__1577 (
            .O(N__14927),
            .I(N__14891));
    LocalMux I__1576 (
            .O(N__14922),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__1575 (
            .O(N__14919),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1574 (
            .O(N__14916),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1573 (
            .O(N__14911),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    LocalMux I__1572 (
            .O(N__14904),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    Odrv4 I__1571 (
            .O(N__14891),
            .I(\this_vga_signals.mult1_un54_sum_axb2_i ));
    InMux I__1570 (
            .O(N__14878),
            .I(N__14875));
    LocalMux I__1569 (
            .O(N__14875),
            .I(\this_vga_signals.g3_0_1 ));
    CascadeMux I__1568 (
            .O(N__14872),
            .I(N__14869));
    InMux I__1567 (
            .O(N__14869),
            .I(N__14866));
    LocalMux I__1566 (
            .O(N__14866),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_c_0 ));
    InMux I__1565 (
            .O(N__14863),
            .I(N__14860));
    LocalMux I__1564 (
            .O(N__14860),
            .I(N__14857));
    Odrv4 I__1563 (
            .O(N__14857),
            .I(\this_vga_signals.mult1_un75_sum_ac0_3_d ));
    InMux I__1562 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__1561 (
            .O(N__14851),
            .I(\this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2 ));
    CascadeMux I__1560 (
            .O(N__14848),
            .I(\this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_ ));
    InMux I__1559 (
            .O(N__14845),
            .I(N__14842));
    LocalMux I__1558 (
            .O(N__14842),
            .I(\this_vga_signals.vaddress_m6_0 ));
    CascadeMux I__1557 (
            .O(N__14839),
            .I(N__14836));
    InMux I__1556 (
            .O(N__14836),
            .I(N__14833));
    LocalMux I__1555 (
            .O(N__14833),
            .I(N__14830));
    Span4Mux_h I__1554 (
            .O(N__14830),
            .I(N__14827));
    Span4Mux_v I__1553 (
            .O(N__14827),
            .I(N__14824));
    Span4Mux_v I__1552 (
            .O(N__14824),
            .I(N__14821));
    Span4Mux_v I__1551 (
            .O(N__14821),
            .I(N__14818));
    Odrv4 I__1550 (
            .O(N__14818),
            .I(M_this_vga_signals_address_7));
    InMux I__1549 (
            .O(N__14815),
            .I(N__14809));
    InMux I__1548 (
            .O(N__14814),
            .I(N__14806));
    InMux I__1547 (
            .O(N__14813),
            .I(N__14803));
    InMux I__1546 (
            .O(N__14812),
            .I(N__14800));
    LocalMux I__1545 (
            .O(N__14809),
            .I(\this_vga_signals.mult1_un61_sum_ac0_4 ));
    LocalMux I__1544 (
            .O(N__14806),
            .I(\this_vga_signals.mult1_un61_sum_ac0_4 ));
    LocalMux I__1543 (
            .O(N__14803),
            .I(\this_vga_signals.mult1_un61_sum_ac0_4 ));
    LocalMux I__1542 (
            .O(N__14800),
            .I(\this_vga_signals.mult1_un61_sum_ac0_4 ));
    InMux I__1541 (
            .O(N__14791),
            .I(N__14788));
    LocalMux I__1540 (
            .O(N__14788),
            .I(N__14785));
    Odrv12 I__1539 (
            .O(N__14785),
            .I(\this_vga_signals.g0_0 ));
    CascadeMux I__1538 (
            .O(N__14782),
            .I(N__14779));
    InMux I__1537 (
            .O(N__14779),
            .I(N__14776));
    LocalMux I__1536 (
            .O(N__14776),
            .I(\this_vga_signals.g0_0_0_0 ));
    InMux I__1535 (
            .O(N__14773),
            .I(N__14770));
    LocalMux I__1534 (
            .O(N__14770),
            .I(\this_vga_signals.g3 ));
    InMux I__1533 (
            .O(N__14767),
            .I(N__14764));
    LocalMux I__1532 (
            .O(N__14764),
            .I(N__14761));
    Odrv12 I__1531 (
            .O(N__14761),
            .I(\this_vga_signals.g0_0_0_a2_2_0 ));
    InMux I__1530 (
            .O(N__14758),
            .I(N__14755));
    LocalMux I__1529 (
            .O(N__14755),
            .I(\this_vga_signals.g0_6_0_a2_3 ));
    CascadeMux I__1528 (
            .O(N__14752),
            .I(\this_vga_signals.N_12_0_0_cascade_ ));
    InMux I__1527 (
            .O(N__14749),
            .I(N__14745));
    CascadeMux I__1526 (
            .O(N__14748),
            .I(N__14741));
    LocalMux I__1525 (
            .O(N__14745),
            .I(N__14735));
    InMux I__1524 (
            .O(N__14744),
            .I(N__14732));
    InMux I__1523 (
            .O(N__14741),
            .I(N__14729));
    InMux I__1522 (
            .O(N__14740),
            .I(N__14722));
    InMux I__1521 (
            .O(N__14739),
            .I(N__14722));
    InMux I__1520 (
            .O(N__14738),
            .I(N__14722));
    Odrv4 I__1519 (
            .O(N__14735),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1518 (
            .O(N__14732),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1517 (
            .O(N__14729),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    LocalMux I__1516 (
            .O(N__14722),
            .I(\this_vga_signals.mult1_un68_sum_c3 ));
    InMux I__1515 (
            .O(N__14713),
            .I(N__14710));
    LocalMux I__1514 (
            .O(N__14710),
            .I(\this_vga_signals.g0_1_1 ));
    InMux I__1513 (
            .O(N__14707),
            .I(N__14700));
    InMux I__1512 (
            .O(N__14706),
            .I(N__14700));
    InMux I__1511 (
            .O(N__14705),
            .I(N__14697));
    LocalMux I__1510 (
            .O(N__14700),
            .I(N__14687));
    LocalMux I__1509 (
            .O(N__14697),
            .I(N__14684));
    InMux I__1508 (
            .O(N__14696),
            .I(N__14681));
    InMux I__1507 (
            .O(N__14695),
            .I(N__14678));
    InMux I__1506 (
            .O(N__14694),
            .I(N__14675));
    InMux I__1505 (
            .O(N__14693),
            .I(N__14672));
    InMux I__1504 (
            .O(N__14692),
            .I(N__14667));
    InMux I__1503 (
            .O(N__14691),
            .I(N__14667));
    InMux I__1502 (
            .O(N__14690),
            .I(N__14664));
    Odrv4 I__1501 (
            .O(N__14687),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__1500 (
            .O(N__14684),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1499 (
            .O(N__14681),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1498 (
            .O(N__14678),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1497 (
            .O(N__14675),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1496 (
            .O(N__14672),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1495 (
            .O(N__14667),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__1494 (
            .O(N__14664),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    InMux I__1493 (
            .O(N__14647),
            .I(N__14644));
    LocalMux I__1492 (
            .O(N__14644),
            .I(\this_vga_signals.g0_0_i_a5_1 ));
    InMux I__1491 (
            .O(N__14641),
            .I(N__14638));
    LocalMux I__1490 (
            .O(N__14638),
            .I(N__14635));
    Span4Mux_v I__1489 (
            .O(N__14635),
            .I(N__14632));
    Odrv4 I__1488 (
            .O(N__14632),
            .I(\this_vga_signals.N_8 ));
    CascadeMux I__1487 (
            .O(N__14629),
            .I(\this_vga_signals.N_6_0_cascade_ ));
    InMux I__1486 (
            .O(N__14626),
            .I(N__14623));
    LocalMux I__1485 (
            .O(N__14623),
            .I(\this_vga_signals.g0_1 ));
    InMux I__1484 (
            .O(N__14620),
            .I(N__14617));
    LocalMux I__1483 (
            .O(N__14617),
            .I(\this_vga_signals.g3_0_0 ));
    InMux I__1482 (
            .O(N__14614),
            .I(N__14611));
    LocalMux I__1481 (
            .O(N__14611),
            .I(\this_vga_signals.g3_1_0 ));
    CascadeMux I__1480 (
            .O(N__14608),
            .I(N__14605));
    InMux I__1479 (
            .O(N__14605),
            .I(N__14602));
    LocalMux I__1478 (
            .O(N__14602),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_0 ));
    InMux I__1477 (
            .O(N__14599),
            .I(N__14596));
    LocalMux I__1476 (
            .O(N__14596),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_0_2 ));
    InMux I__1475 (
            .O(N__14593),
            .I(N__14587));
    InMux I__1474 (
            .O(N__14592),
            .I(N__14584));
    InMux I__1473 (
            .O(N__14591),
            .I(N__14577));
    InMux I__1472 (
            .O(N__14590),
            .I(N__14577));
    LocalMux I__1471 (
            .O(N__14587),
            .I(N__14574));
    LocalMux I__1470 (
            .O(N__14584),
            .I(N__14571));
    InMux I__1469 (
            .O(N__14583),
            .I(N__14562));
    InMux I__1468 (
            .O(N__14582),
            .I(N__14559));
    LocalMux I__1467 (
            .O(N__14577),
            .I(N__14552));
    Span4Mux_v I__1466 (
            .O(N__14574),
            .I(N__14552));
    Span4Mux_s2_h I__1465 (
            .O(N__14571),
            .I(N__14552));
    InMux I__1464 (
            .O(N__14570),
            .I(N__14549));
    InMux I__1463 (
            .O(N__14569),
            .I(N__14544));
    InMux I__1462 (
            .O(N__14568),
            .I(N__14544));
    InMux I__1461 (
            .O(N__14567),
            .I(N__14537));
    InMux I__1460 (
            .O(N__14566),
            .I(N__14537));
    InMux I__1459 (
            .O(N__14565),
            .I(N__14537));
    LocalMux I__1458 (
            .O(N__14562),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1457 (
            .O(N__14559),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    Odrv4 I__1456 (
            .O(N__14552),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1455 (
            .O(N__14549),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1454 (
            .O(N__14544),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    LocalMux I__1453 (
            .O(N__14537),
            .I(\this_vga_signals.mult1_un40_sum_axb1_i ));
    InMux I__1452 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__1451 (
            .O(N__14521),
            .I(N__14518));
    Odrv4 I__1450 (
            .O(N__14518),
            .I(\this_vga_signals.g0_15 ));
    CascadeMux I__1449 (
            .O(N__14515),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_ ));
    CascadeMux I__1448 (
            .O(N__14512),
            .I(\this_vga_signals.N_1_4_1_cascade_ ));
    CascadeMux I__1447 (
            .O(N__14509),
            .I(\this_vga_signals.mult1_un40_sum_c2_1_cascade_ ));
    CascadeMux I__1446 (
            .O(N__14506),
            .I(\this_vga_signals.mult1_un40_sum_c2_0_cascade_ ));
    CascadeMux I__1445 (
            .O(N__14503),
            .I(\this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_ ));
    InMux I__1444 (
            .O(N__14500),
            .I(N__14497));
    LocalMux I__1443 (
            .O(N__14497),
            .I(\this_vga_signals.mult1_un40_sum_c2_2 ));
    InMux I__1442 (
            .O(N__14494),
            .I(N__14491));
    LocalMux I__1441 (
            .O(N__14491),
            .I(N__14488));
    Odrv4 I__1440 (
            .O(N__14488),
            .I(\this_vga_signals.N_4_3 ));
    InMux I__1439 (
            .O(N__14485),
            .I(N__14482));
    LocalMux I__1438 (
            .O(N__14482),
            .I(\this_vga_signals.g1_1_1 ));
    InMux I__1437 (
            .O(N__14479),
            .I(N__14476));
    LocalMux I__1436 (
            .O(N__14476),
            .I(\this_vga_signals.mult1_un40_sum_ac0_2 ));
    InMux I__1435 (
            .O(N__14473),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    CascadeMux I__1434 (
            .O(N__14470),
            .I(N__14467));
    InMux I__1433 (
            .O(N__14467),
            .I(N__14464));
    LocalMux I__1432 (
            .O(N__14464),
            .I(N__14461));
    Odrv4 I__1431 (
            .O(N__14461),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1 ));
    InMux I__1430 (
            .O(N__14458),
            .I(N__14455));
    LocalMux I__1429 (
            .O(N__14455),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2_2 ));
    InMux I__1428 (
            .O(N__14452),
            .I(N__14447));
    InMux I__1427 (
            .O(N__14451),
            .I(N__14444));
    InMux I__1426 (
            .O(N__14450),
            .I(N__14441));
    LocalMux I__1425 (
            .O(N__14447),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__1424 (
            .O(N__14444),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    LocalMux I__1423 (
            .O(N__14441),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    InMux I__1422 (
            .O(N__14434),
            .I(N__14431));
    LocalMux I__1421 (
            .O(N__14431),
            .I(N__14427));
    InMux I__1420 (
            .O(N__14430),
            .I(N__14424));
    Odrv4 I__1419 (
            .O(N__14427),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__1418 (
            .O(N__14424),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__1417 (
            .O(N__14419),
            .I(N__14416));
    LocalMux I__1416 (
            .O(N__14416),
            .I(N__14410));
    InMux I__1415 (
            .O(N__14415),
            .I(N__14405));
    InMux I__1414 (
            .O(N__14414),
            .I(N__14405));
    InMux I__1413 (
            .O(N__14413),
            .I(N__14402));
    Odrv4 I__1412 (
            .O(N__14410),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__1411 (
            .O(N__14405),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__1410 (
            .O(N__14402),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    InMux I__1409 (
            .O(N__14395),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__1408 (
            .O(N__14392),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__1407 (
            .O(N__14389),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__1406 (
            .O(N__14386),
            .I(N__14383));
    LocalMux I__1405 (
            .O(N__14383),
            .I(N__14379));
    InMux I__1404 (
            .O(N__14382),
            .I(N__14376));
    Span4Mux_s2_h I__1403 (
            .O(N__14379),
            .I(N__14372));
    LocalMux I__1402 (
            .O(N__14376),
            .I(N__14369));
    InMux I__1401 (
            .O(N__14375),
            .I(N__14366));
    Odrv4 I__1400 (
            .O(N__14372),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__1399 (
            .O(N__14369),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    LocalMux I__1398 (
            .O(N__14366),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__1397 (
            .O(N__14359),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__1396 (
            .O(N__14356),
            .I(N__14350));
    InMux I__1395 (
            .O(N__14355),
            .I(N__14350));
    LocalMux I__1394 (
            .O(N__14350),
            .I(N__14347));
    Span4Mux_v I__1393 (
            .O(N__14347),
            .I(N__14343));
    InMux I__1392 (
            .O(N__14346),
            .I(N__14340));
    Odrv4 I__1391 (
            .O(N__14343),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    LocalMux I__1390 (
            .O(N__14340),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__1389 (
            .O(N__14335),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__1388 (
            .O(N__14332),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__1387 (
            .O(N__14329),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__1386 (
            .O(N__14326),
            .I(bfn_3_10_0_));
    CascadeMux I__1385 (
            .O(N__14323),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ));
    InMux I__1384 (
            .O(N__14320),
            .I(N__14317));
    LocalMux I__1383 (
            .O(N__14317),
            .I(\this_vga_signals.g0_2 ));
    CascadeMux I__1382 (
            .O(N__14314),
            .I(\this_vga_signals.mult1_un68_sum_0_3_cascade_ ));
    InMux I__1381 (
            .O(N__14311),
            .I(N__14308));
    LocalMux I__1380 (
            .O(N__14308),
            .I(\this_vga_signals.mult1_un75_sum_ac0_1 ));
    InMux I__1379 (
            .O(N__14305),
            .I(N__14294));
    InMux I__1378 (
            .O(N__14304),
            .I(N__14294));
    InMux I__1377 (
            .O(N__14303),
            .I(N__14294));
    CascadeMux I__1376 (
            .O(N__14302),
            .I(N__14289));
    CascadeMux I__1375 (
            .O(N__14301),
            .I(N__14286));
    LocalMux I__1374 (
            .O(N__14294),
            .I(N__14278));
    InMux I__1373 (
            .O(N__14293),
            .I(N__14273));
    InMux I__1372 (
            .O(N__14292),
            .I(N__14273));
    InMux I__1371 (
            .O(N__14289),
            .I(N__14270));
    InMux I__1370 (
            .O(N__14286),
            .I(N__14267));
    InMux I__1369 (
            .O(N__14285),
            .I(N__14259));
    InMux I__1368 (
            .O(N__14284),
            .I(N__14259));
    InMux I__1367 (
            .O(N__14283),
            .I(N__14252));
    InMux I__1366 (
            .O(N__14282),
            .I(N__14252));
    InMux I__1365 (
            .O(N__14281),
            .I(N__14252));
    Span4Mux_v I__1364 (
            .O(N__14278),
            .I(N__14243));
    LocalMux I__1363 (
            .O(N__14273),
            .I(N__14243));
    LocalMux I__1362 (
            .O(N__14270),
            .I(N__14243));
    LocalMux I__1361 (
            .O(N__14267),
            .I(N__14243));
    InMux I__1360 (
            .O(N__14266),
            .I(N__14236));
    InMux I__1359 (
            .O(N__14265),
            .I(N__14236));
    InMux I__1358 (
            .O(N__14264),
            .I(N__14236));
    LocalMux I__1357 (
            .O(N__14259),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1356 (
            .O(N__14252),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    Odrv4 I__1355 (
            .O(N__14243),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    LocalMux I__1354 (
            .O(N__14236),
            .I(\this_vga_signals.mult1_un47_sum_c3 ));
    InMux I__1353 (
            .O(N__14227),
            .I(N__14224));
    LocalMux I__1352 (
            .O(N__14224),
            .I(N__14220));
    InMux I__1351 (
            .O(N__14223),
            .I(N__14214));
    Span4Mux_h I__1350 (
            .O(N__14220),
            .I(N__14211));
    InMux I__1349 (
            .O(N__14219),
            .I(N__14204));
    InMux I__1348 (
            .O(N__14218),
            .I(N__14204));
    InMux I__1347 (
            .O(N__14217),
            .I(N__14204));
    LocalMux I__1346 (
            .O(N__14214),
            .I(N__14201));
    Odrv4 I__1345 (
            .O(N__14211),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    LocalMux I__1344 (
            .O(N__14204),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    Odrv4 I__1343 (
            .O(N__14201),
            .I(\this_vga_signals.mult1_un61_sum_c2_0 ));
    CascadeMux I__1342 (
            .O(N__14194),
            .I(\this_vga_signals.g3_0_a2_2_cascade_ ));
    InMux I__1341 (
            .O(N__14191),
            .I(N__14184));
    InMux I__1340 (
            .O(N__14190),
            .I(N__14184));
    InMux I__1339 (
            .O(N__14189),
            .I(N__14181));
    LocalMux I__1338 (
            .O(N__14184),
            .I(\this_vga_signals.mult1_un75_sum_axb2 ));
    LocalMux I__1337 (
            .O(N__14181),
            .I(\this_vga_signals.mult1_un75_sum_axb2 ));
    InMux I__1336 (
            .O(N__14176),
            .I(N__14173));
    LocalMux I__1335 (
            .O(N__14173),
            .I(\this_vga_signals.g0_1_0 ));
    InMux I__1334 (
            .O(N__14170),
            .I(N__14166));
    InMux I__1333 (
            .O(N__14169),
            .I(N__14163));
    LocalMux I__1332 (
            .O(N__14166),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    LocalMux I__1331 (
            .O(N__14163),
            .I(\this_vga_signals.mult1_un61_sum_c3_0 ));
    InMux I__1330 (
            .O(N__14158),
            .I(N__14155));
    LocalMux I__1329 (
            .O(N__14155),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0 ));
    InMux I__1328 (
            .O(N__14152),
            .I(N__14149));
    LocalMux I__1327 (
            .O(N__14149),
            .I(\this_vga_signals.if_i4_mux_0 ));
    CascadeMux I__1326 (
            .O(N__14146),
            .I(\this_vga_signals.vaddress_N_3_i_0_0_cascade_ ));
    InMux I__1325 (
            .O(N__14143),
            .I(N__14140));
    LocalMux I__1324 (
            .O(N__14140),
            .I(N__14137));
    Odrv4 I__1323 (
            .O(N__14137),
            .I(\this_vga_signals.g2_4_0 ));
    CascadeMux I__1322 (
            .O(N__14134),
            .I(N__14131));
    InMux I__1321 (
            .O(N__14131),
            .I(N__14128));
    LocalMux I__1320 (
            .O(N__14128),
            .I(\this_vga_signals.g2_0_0 ));
    InMux I__1319 (
            .O(N__14125),
            .I(N__14122));
    LocalMux I__1318 (
            .O(N__14122),
            .I(\this_vga_signals.g0_4_0 ));
    InMux I__1317 (
            .O(N__14119),
            .I(N__14115));
    InMux I__1316 (
            .O(N__14118),
            .I(N__14112));
    LocalMux I__1315 (
            .O(N__14115),
            .I(N__14109));
    LocalMux I__1314 (
            .O(N__14112),
            .I(N__14106));
    Span4Mux_v I__1313 (
            .O(N__14109),
            .I(N__14103));
    Odrv12 I__1312 (
            .O(N__14106),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0 ));
    Odrv4 I__1311 (
            .O(N__14103),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0 ));
    InMux I__1310 (
            .O(N__14098),
            .I(N__14095));
    LocalMux I__1309 (
            .O(N__14095),
            .I(N__14092));
    Odrv4 I__1308 (
            .O(N__14092),
            .I(\this_vga_signals.g0_0_6 ));
    InMux I__1307 (
            .O(N__14089),
            .I(N__14086));
    LocalMux I__1306 (
            .O(N__14086),
            .I(\this_vga_signals.g1_0_0_0_0 ));
    CascadeMux I__1305 (
            .O(N__14083),
            .I(N__14079));
    CascadeMux I__1304 (
            .O(N__14082),
            .I(N__14076));
    InMux I__1303 (
            .O(N__14079),
            .I(N__14072));
    InMux I__1302 (
            .O(N__14076),
            .I(N__14069));
    InMux I__1301 (
            .O(N__14075),
            .I(N__14066));
    LocalMux I__1300 (
            .O(N__14072),
            .I(N__14056));
    LocalMux I__1299 (
            .O(N__14069),
            .I(N__14056));
    LocalMux I__1298 (
            .O(N__14066),
            .I(N__14053));
    InMux I__1297 (
            .O(N__14065),
            .I(N__14046));
    InMux I__1296 (
            .O(N__14064),
            .I(N__14046));
    InMux I__1295 (
            .O(N__14063),
            .I(N__14046));
    InMux I__1294 (
            .O(N__14062),
            .I(N__14041));
    InMux I__1293 (
            .O(N__14061),
            .I(N__14041));
    Odrv4 I__1292 (
            .O(N__14056),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4 ));
    Odrv4 I__1291 (
            .O(N__14053),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4 ));
    LocalMux I__1290 (
            .O(N__14046),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4 ));
    LocalMux I__1289 (
            .O(N__14041),
            .I(\this_vga_signals.mult1_un54_sum_ac0_4 ));
    InMux I__1288 (
            .O(N__14032),
            .I(N__14029));
    LocalMux I__1287 (
            .O(N__14029),
            .I(N__14026));
    Span4Mux_v I__1286 (
            .O(N__14026),
            .I(N__14023));
    Odrv4 I__1285 (
            .O(N__14023),
            .I(\this_vga_signals.g3_0 ));
    InMux I__1284 (
            .O(N__14020),
            .I(N__14017));
    LocalMux I__1283 (
            .O(N__14017),
            .I(\this_vga_signals.N_3_2 ));
    InMux I__1282 (
            .O(N__14014),
            .I(N__14008));
    InMux I__1281 (
            .O(N__14013),
            .I(N__14005));
    InMux I__1280 (
            .O(N__14012),
            .I(N__14000));
    InMux I__1279 (
            .O(N__14011),
            .I(N__14000));
    LocalMux I__1278 (
            .O(N__14008),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__1277 (
            .O(N__14005),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    LocalMux I__1276 (
            .O(N__14000),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1 ));
    CascadeMux I__1275 (
            .O(N__13993),
            .I(N__13987));
    InMux I__1274 (
            .O(N__13992),
            .I(N__13977));
    InMux I__1273 (
            .O(N__13991),
            .I(N__13977));
    InMux I__1272 (
            .O(N__13990),
            .I(N__13977));
    InMux I__1271 (
            .O(N__13987),
            .I(N__13964));
    InMux I__1270 (
            .O(N__13986),
            .I(N__13961));
    InMux I__1269 (
            .O(N__13985),
            .I(N__13956));
    InMux I__1268 (
            .O(N__13984),
            .I(N__13956));
    LocalMux I__1267 (
            .O(N__13977),
            .I(N__13953));
    InMux I__1266 (
            .O(N__13976),
            .I(N__13944));
    InMux I__1265 (
            .O(N__13975),
            .I(N__13944));
    InMux I__1264 (
            .O(N__13974),
            .I(N__13944));
    InMux I__1263 (
            .O(N__13973),
            .I(N__13944));
    InMux I__1262 (
            .O(N__13972),
            .I(N__13935));
    InMux I__1261 (
            .O(N__13971),
            .I(N__13935));
    InMux I__1260 (
            .O(N__13970),
            .I(N__13935));
    InMux I__1259 (
            .O(N__13969),
            .I(N__13935));
    InMux I__1258 (
            .O(N__13968),
            .I(N__13930));
    InMux I__1257 (
            .O(N__13967),
            .I(N__13930));
    LocalMux I__1256 (
            .O(N__13964),
            .I(N__13927));
    LocalMux I__1255 (
            .O(N__13961),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1254 (
            .O(N__13956),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__1253 (
            .O(N__13953),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1252 (
            .O(N__13944),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1251 (
            .O(N__13935),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__1250 (
            .O(N__13930),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv12 I__1249 (
            .O(N__13927),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__1248 (
            .O(N__13912),
            .I(N__13909));
    LocalMux I__1247 (
            .O(N__13909),
            .I(\this_vga_signals.g2_0_0_0 ));
    InMux I__1246 (
            .O(N__13906),
            .I(N__13903));
    LocalMux I__1245 (
            .O(N__13903),
            .I(\this_vga_signals.g3_x0 ));
    InMux I__1244 (
            .O(N__13900),
            .I(N__13893));
    InMux I__1243 (
            .O(N__13899),
            .I(N__13893));
    CascadeMux I__1242 (
            .O(N__13898),
            .I(N__13888));
    LocalMux I__1241 (
            .O(N__13893),
            .I(N__13882));
    InMux I__1240 (
            .O(N__13892),
            .I(N__13877));
    InMux I__1239 (
            .O(N__13891),
            .I(N__13877));
    InMux I__1238 (
            .O(N__13888),
            .I(N__13868));
    InMux I__1237 (
            .O(N__13887),
            .I(N__13868));
    InMux I__1236 (
            .O(N__13886),
            .I(N__13868));
    InMux I__1235 (
            .O(N__13885),
            .I(N__13868));
    Odrv4 I__1234 (
            .O(N__13882),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1233 (
            .O(N__13877),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    LocalMux I__1232 (
            .O(N__13868),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    InMux I__1231 (
            .O(N__13861),
            .I(N__13858));
    LocalMux I__1230 (
            .O(N__13858),
            .I(\this_vga_signals.g3_x1 ));
    InMux I__1229 (
            .O(N__13855),
            .I(N__13846));
    InMux I__1228 (
            .O(N__13854),
            .I(N__13846));
    InMux I__1227 (
            .O(N__13853),
            .I(N__13843));
    InMux I__1226 (
            .O(N__13852),
            .I(N__13840));
    InMux I__1225 (
            .O(N__13851),
            .I(N__13837));
    LocalMux I__1224 (
            .O(N__13846),
            .I(N__13834));
    LocalMux I__1223 (
            .O(N__13843),
            .I(N__13831));
    LocalMux I__1222 (
            .O(N__13840),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    LocalMux I__1221 (
            .O(N__13837),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    Odrv4 I__1220 (
            .O(N__13834),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    Odrv4 I__1219 (
            .O(N__13831),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i ));
    CascadeMux I__1218 (
            .O(N__13822),
            .I(N__13819));
    InMux I__1217 (
            .O(N__13819),
            .I(N__13816));
    LocalMux I__1216 (
            .O(N__13816),
            .I(\this_vga_signals.mult1_un61_sum_ac0_1 ));
    InMux I__1215 (
            .O(N__13813),
            .I(N__13810));
    LocalMux I__1214 (
            .O(N__13810),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_3 ));
    CascadeMux I__1213 (
            .O(N__13807),
            .I(\this_vga_signals.g1_0_0_2_cascade_ ));
    CascadeMux I__1212 (
            .O(N__13804),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__1211 (
            .O(N__13801),
            .I(N__13798));
    LocalMux I__1210 (
            .O(N__13798),
            .I(\this_vga_signals.g0_0_0_1_0 ));
    CascadeMux I__1209 (
            .O(N__13795),
            .I(N__13788));
    InMux I__1208 (
            .O(N__13794),
            .I(N__13783));
    InMux I__1207 (
            .O(N__13793),
            .I(N__13783));
    InMux I__1206 (
            .O(N__13792),
            .I(N__13780));
    InMux I__1205 (
            .O(N__13791),
            .I(N__13777));
    InMux I__1204 (
            .O(N__13788),
            .I(N__13774));
    LocalMux I__1203 (
            .O(N__13783),
            .I(N__13771));
    LocalMux I__1202 (
            .O(N__13780),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__1201 (
            .O(N__13777),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__1200 (
            .O(N__13774),
            .I(\this_vga_signals.vaddress_6 ));
    Odrv4 I__1199 (
            .O(N__13771),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__1198 (
            .O(N__13762),
            .I(N__13759));
    LocalMux I__1197 (
            .O(N__13759),
            .I(N__13756));
    Odrv4 I__1196 (
            .O(N__13756),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_0 ));
    CascadeMux I__1195 (
            .O(N__13753),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ));
    InMux I__1194 (
            .O(N__13750),
            .I(N__13741));
    InMux I__1193 (
            .O(N__13749),
            .I(N__13741));
    CascadeMux I__1192 (
            .O(N__13748),
            .I(N__13738));
    InMux I__1191 (
            .O(N__13747),
            .I(N__13735));
    InMux I__1190 (
            .O(N__13746),
            .I(N__13732));
    LocalMux I__1189 (
            .O(N__13741),
            .I(N__13729));
    InMux I__1188 (
            .O(N__13738),
            .I(N__13726));
    LocalMux I__1187 (
            .O(N__13735),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    LocalMux I__1186 (
            .O(N__13732),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    Odrv4 I__1185 (
            .O(N__13729),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    LocalMux I__1184 (
            .O(N__13726),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1 ));
    CascadeMux I__1183 (
            .O(N__13717),
            .I(N__13712));
    InMux I__1182 (
            .O(N__13716),
            .I(N__13698));
    InMux I__1181 (
            .O(N__13715),
            .I(N__13698));
    InMux I__1180 (
            .O(N__13712),
            .I(N__13693));
    InMux I__1179 (
            .O(N__13711),
            .I(N__13693));
    InMux I__1178 (
            .O(N__13710),
            .I(N__13688));
    InMux I__1177 (
            .O(N__13709),
            .I(N__13688));
    InMux I__1176 (
            .O(N__13708),
            .I(N__13679));
    InMux I__1175 (
            .O(N__13707),
            .I(N__13679));
    InMux I__1174 (
            .O(N__13706),
            .I(N__13679));
    InMux I__1173 (
            .O(N__13705),
            .I(N__13679));
    InMux I__1172 (
            .O(N__13704),
            .I(N__13674));
    InMux I__1171 (
            .O(N__13703),
            .I(N__13674));
    LocalMux I__1170 (
            .O(N__13698),
            .I(N__13669));
    LocalMux I__1169 (
            .O(N__13693),
            .I(N__13669));
    LocalMux I__1168 (
            .O(N__13688),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__1167 (
            .O(N__13679),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    LocalMux I__1166 (
            .O(N__13674),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    Odrv4 I__1165 (
            .O(N__13669),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2 ));
    CascadeMux I__1164 (
            .O(N__13660),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_4_cascade_ ));
    InMux I__1163 (
            .O(N__13657),
            .I(N__13654));
    LocalMux I__1162 (
            .O(N__13654),
            .I(N__13650));
    InMux I__1161 (
            .O(N__13653),
            .I(N__13647));
    Span4Mux_h I__1160 (
            .O(N__13650),
            .I(N__13644));
    LocalMux I__1159 (
            .O(N__13647),
            .I(\this_vga_signals.g2_1_0 ));
    Odrv4 I__1158 (
            .O(N__13644),
            .I(\this_vga_signals.g2_1_0 ));
    InMux I__1157 (
            .O(N__13639),
            .I(N__13636));
    LocalMux I__1156 (
            .O(N__13636),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2_mb_sn ));
    CascadeMux I__1155 (
            .O(N__13633),
            .I(N__13629));
    InMux I__1154 (
            .O(N__13632),
            .I(N__13625));
    InMux I__1153 (
            .O(N__13629),
            .I(N__13620));
    InMux I__1152 (
            .O(N__13628),
            .I(N__13620));
    LocalMux I__1151 (
            .O(N__13625),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0 ));
    LocalMux I__1150 (
            .O(N__13620),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0 ));
    CascadeMux I__1149 (
            .O(N__13615),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ));
    InMux I__1148 (
            .O(N__13612),
            .I(N__13609));
    LocalMux I__1147 (
            .O(N__13609),
            .I(N__13606));
    Span4Mux_v I__1146 (
            .O(N__13606),
            .I(N__13603));
    Odrv4 I__1145 (
            .O(N__13603),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_1 ));
    CascadeMux I__1144 (
            .O(N__13600),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_ ));
    CascadeMux I__1143 (
            .O(N__13597),
            .I(N__13593));
    InMux I__1142 (
            .O(N__13596),
            .I(N__13590));
    InMux I__1141 (
            .O(N__13593),
            .I(N__13587));
    LocalMux I__1140 (
            .O(N__13590),
            .I(N__13584));
    LocalMux I__1139 (
            .O(N__13587),
            .I(\this_vga_signals.SUM_2_i_i_1_1_3 ));
    Odrv4 I__1138 (
            .O(N__13584),
            .I(\this_vga_signals.SUM_2_i_i_1_1_3 ));
    CascadeMux I__1137 (
            .O(N__13579),
            .I(N__13576));
    InMux I__1136 (
            .O(N__13576),
            .I(N__13573));
    LocalMux I__1135 (
            .O(N__13573),
            .I(\this_vga_signals.mult1_un40_sum_axb1_x0 ));
    InMux I__1134 (
            .O(N__13570),
            .I(N__13567));
    LocalMux I__1133 (
            .O(N__13567),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0 ));
    CascadeMux I__1132 (
            .O(N__13564),
            .I(N__13560));
    InMux I__1131 (
            .O(N__13563),
            .I(N__13557));
    InMux I__1130 (
            .O(N__13560),
            .I(N__13554));
    LocalMux I__1129 (
            .O(N__13557),
            .I(\this_vga_signals.SUM_2_i_i_1_0_3 ));
    LocalMux I__1128 (
            .O(N__13554),
            .I(\this_vga_signals.SUM_2_i_i_1_0_3 ));
    InMux I__1127 (
            .O(N__13549),
            .I(N__13546));
    LocalMux I__1126 (
            .O(N__13546),
            .I(\this_vga_signals.mult1_un40_sum_axb1_x1 ));
    InMux I__1125 (
            .O(N__13543),
            .I(N__13538));
    CascadeMux I__1124 (
            .O(N__13542),
            .I(N__13535));
    CascadeMux I__1123 (
            .O(N__13541),
            .I(N__13531));
    LocalMux I__1122 (
            .O(N__13538),
            .I(N__13528));
    InMux I__1121 (
            .O(N__13535),
            .I(N__13525));
    InMux I__1120 (
            .O(N__13534),
            .I(N__13520));
    InMux I__1119 (
            .O(N__13531),
            .I(N__13520));
    Odrv4 I__1118 (
            .O(N__13528),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1117 (
            .O(N__13525),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    LocalMux I__1116 (
            .O(N__13520),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__1115 (
            .O(N__13513),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_ ));
    InMux I__1114 (
            .O(N__13510),
            .I(N__13507));
    LocalMux I__1113 (
            .O(N__13507),
            .I(N__13501));
    InMux I__1112 (
            .O(N__13506),
            .I(N__13498));
    InMux I__1111 (
            .O(N__13505),
            .I(N__13493));
    InMux I__1110 (
            .O(N__13504),
            .I(N__13493));
    Odrv4 I__1109 (
            .O(N__13501),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1108 (
            .O(N__13498),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    LocalMux I__1107 (
            .O(N__13493),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__1106 (
            .O(N__13486),
            .I(N__13483));
    LocalMux I__1105 (
            .O(N__13483),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns ));
    CascadeMux I__1104 (
            .O(N__13480),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_ ));
    InMux I__1103 (
            .O(N__13477),
            .I(N__13474));
    LocalMux I__1102 (
            .O(N__13474),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2 ));
    CascadeMux I__1101 (
            .O(N__13471),
            .I(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ));
    CascadeMux I__1100 (
            .O(N__13468),
            .I(N__13464));
    CascadeMux I__1099 (
            .O(N__13467),
            .I(N__13461));
    InMux I__1098 (
            .O(N__13464),
            .I(N__13458));
    InMux I__1097 (
            .O(N__13461),
            .I(N__13455));
    LocalMux I__1096 (
            .O(N__13458),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    LocalMux I__1095 (
            .O(N__13455),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    CascadeMux I__1094 (
            .O(N__13450),
            .I(\this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ));
    InMux I__1093 (
            .O(N__13447),
            .I(N__13442));
    InMux I__1092 (
            .O(N__13446),
            .I(N__13437));
    InMux I__1091 (
            .O(N__13445),
            .I(N__13437));
    LocalMux I__1090 (
            .O(N__13442),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__1089 (
            .O(N__13437),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    CascadeMux I__1088 (
            .O(N__13432),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_ ));
    InMux I__1087 (
            .O(N__13429),
            .I(N__13426));
    LocalMux I__1086 (
            .O(N__13426),
            .I(\this_vga_signals.g1_0_0_1 ));
    IoInMux I__1085 (
            .O(N__13423),
            .I(N__13420));
    LocalMux I__1084 (
            .O(N__13420),
            .I(N__13417));
    Span4Mux_s2_h I__1083 (
            .O(N__13417),
            .I(N__13414));
    Span4Mux_v I__1082 (
            .O(N__13414),
            .I(N__13411));
    Odrv4 I__1081 (
            .O(N__13411),
            .I(port_data_rw_0_i));
    CascadeMux I__1080 (
            .O(N__13408),
            .I(N__13405));
    InMux I__1079 (
            .O(N__13405),
            .I(N__13402));
    LocalMux I__1078 (
            .O(N__13402),
            .I(\this_vga_signals.g2_2_0 ));
    IoInMux I__1077 (
            .O(N__13399),
            .I(N__13396));
    LocalMux I__1076 (
            .O(N__13396),
            .I(N__13393));
    Span4Mux_s2_h I__1075 (
            .O(N__13393),
            .I(N__13390));
    Odrv4 I__1074 (
            .O(N__13390),
            .I(rgb_c_0));
    IoInMux I__1073 (
            .O(N__13387),
            .I(N__13384));
    LocalMux I__1072 (
            .O(N__13384),
            .I(N__13381));
    Span4Mux_s1_h I__1071 (
            .O(N__13381),
            .I(N__13378));
    Span4Mux_v I__1070 (
            .O(N__13378),
            .I(N__13375));
    Span4Mux_v I__1069 (
            .O(N__13375),
            .I(N__13372));
    Odrv4 I__1068 (
            .O(N__13372),
            .I(rgb_c_1));
    CascadeMux I__1067 (
            .O(N__13369),
            .I(N__13366));
    InMux I__1066 (
            .O(N__13366),
            .I(N__13363));
    LocalMux I__1065 (
            .O(N__13363),
            .I(N__13360));
    Odrv4 I__1064 (
            .O(N__13360),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_2 ));
    CascadeMux I__1063 (
            .O(N__13357),
            .I(N__13354));
    InMux I__1062 (
            .O(N__13354),
            .I(N__13351));
    LocalMux I__1061 (
            .O(N__13351),
            .I(N__13348));
    Odrv4 I__1060 (
            .O(N__13348),
            .I(\this_vga_signals.g1_1_0 ));
    CascadeMux I__1059 (
            .O(N__13345),
            .I(\this_vga_signals.g1_4_cascade_ ));
    IoInMux I__1058 (
            .O(N__13342),
            .I(N__13339));
    LocalMux I__1057 (
            .O(N__13339),
            .I(N__13336));
    Span12Mux_s0_h I__1056 (
            .O(N__13336),
            .I(N__13333));
    Span12Mux_v I__1055 (
            .O(N__13333),
            .I(N__13330));
    Odrv12 I__1054 (
            .O(N__13330),
            .I(rgb_c_4));
    InMux I__1053 (
            .O(N__13327),
            .I(N__13322));
    InMux I__1052 (
            .O(N__13326),
            .I(N__13317));
    InMux I__1051 (
            .O(N__13325),
            .I(N__13317));
    LocalMux I__1050 (
            .O(N__13322),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    LocalMux I__1049 (
            .O(N__13317),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_1 ));
    InMux I__1048 (
            .O(N__13312),
            .I(N__13309));
    LocalMux I__1047 (
            .O(N__13309),
            .I(N__13306));
    Odrv4 I__1046 (
            .O(N__13306),
            .I(\this_vga_signals.vaddress_m2_2 ));
    InMux I__1045 (
            .O(N__13303),
            .I(N__13300));
    LocalMux I__1044 (
            .O(N__13300),
            .I(N__13297));
    IoSpan4Mux I__1043 (
            .O(N__13297),
            .I(N__13294));
    Odrv4 I__1042 (
            .O(N__13294),
            .I(port_clk_c));
    InMux I__1041 (
            .O(N__13291),
            .I(N__13288));
    LocalMux I__1040 (
            .O(N__13288),
            .I(N__13285));
    Odrv12 I__1039 (
            .O(N__13285),
            .I(\this_vga_signals.g2 ));
    InMux I__1038 (
            .O(N__13282),
            .I(N__13279));
    LocalMux I__1037 (
            .O(N__13279),
            .I(N__13275));
    InMux I__1036 (
            .O(N__13278),
            .I(N__13272));
    Span4Mux_v I__1035 (
            .O(N__13275),
            .I(N__13267));
    LocalMux I__1034 (
            .O(N__13272),
            .I(N__13267));
    Odrv4 I__1033 (
            .O(N__13267),
            .I(\this_vga_signals.g1 ));
    IoInMux I__1032 (
            .O(N__13264),
            .I(N__13261));
    LocalMux I__1031 (
            .O(N__13261),
            .I(\this_vga_signals.N_935_0 ));
    InMux I__1030 (
            .O(N__13258),
            .I(N__13255));
    LocalMux I__1029 (
            .O(N__13255),
            .I(N__13252));
    Odrv12 I__1028 (
            .O(N__13252),
            .I(\this_vga_signals.g3_2 ));
    CascadeMux I__1027 (
            .O(N__13249),
            .I(\this_vga_signals.mult1_un75_sum_axb1_3_cascade_ ));
    InMux I__1026 (
            .O(N__13246),
            .I(N__13243));
    LocalMux I__1025 (
            .O(N__13243),
            .I(N__13240));
    Span4Mux_v I__1024 (
            .O(N__13240),
            .I(N__13237));
    Odrv4 I__1023 (
            .O(N__13237),
            .I(\this_vga_signals.vaddress_m2_1 ));
    InMux I__1022 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__1021 (
            .O(N__13231),
            .I(N__13228));
    Odrv12 I__1020 (
            .O(N__13228),
            .I(\this_vga_signals.if_N_9_i ));
    InMux I__1019 (
            .O(N__13225),
            .I(N__13222));
    LocalMux I__1018 (
            .O(N__13222),
            .I(\this_vga_signals.if_m1_0 ));
    CascadeMux I__1017 (
            .O(N__13219),
            .I(\this_vga_signals.mult1_un68_sum_c3_cascade_ ));
    InMux I__1016 (
            .O(N__13216),
            .I(N__13213));
    LocalMux I__1015 (
            .O(N__13213),
            .I(N__13210));
    Odrv4 I__1014 (
            .O(N__13210),
            .I(\this_vga_signals.mult1_un61_sum_axb2_i_0 ));
    InMux I__1013 (
            .O(N__13207),
            .I(N__13204));
    LocalMux I__1012 (
            .O(N__13204),
            .I(\this_vga_signals.g2_3 ));
    CascadeMux I__1011 (
            .O(N__13201),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_ ));
    CascadeMux I__1010 (
            .O(N__13198),
            .I(\this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_ ));
    InMux I__1009 (
            .O(N__13195),
            .I(N__13191));
    InMux I__1008 (
            .O(N__13194),
            .I(N__13188));
    LocalMux I__1007 (
            .O(N__13191),
            .I(\this_vga_signals.mult1_un75_sum_axb1_3_1 ));
    LocalMux I__1006 (
            .O(N__13188),
            .I(\this_vga_signals.mult1_un75_sum_axb1_3_1 ));
    CascadeMux I__1005 (
            .O(N__13183),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ));
    CascadeMux I__1004 (
            .O(N__13180),
            .I(\this_vga_signals.g1_0_0_0_cascade_ ));
    InMux I__1003 (
            .O(N__13177),
            .I(N__13174));
    LocalMux I__1002 (
            .O(N__13174),
            .I(\this_vga_signals.g1_0_0_0 ));
    InMux I__1001 (
            .O(N__13171),
            .I(N__13168));
    LocalMux I__1000 (
            .O(N__13168),
            .I(N__13165));
    Odrv12 I__999 (
            .O(N__13165),
            .I(\this_vga_signals.g2_1 ));
    CascadeMux I__998 (
            .O(N__13162),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ));
    CascadeMux I__997 (
            .O(N__13159),
            .I(\this_vga_signals.g2_1_0_cascade_ ));
    CascadeMux I__996 (
            .O(N__13156),
            .I(\this_vga_signals.g2_0_cascade_ ));
    CascadeMux I__995 (
            .O(N__13153),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1_cascade_ ));
    CascadeMux I__994 (
            .O(N__13150),
            .I(N__13147));
    InMux I__993 (
            .O(N__13147),
            .I(N__13144));
    LocalMux I__992 (
            .O(N__13144),
            .I(N__13141));
    Odrv4 I__991 (
            .O(N__13141),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ));
    InMux I__990 (
            .O(N__13138),
            .I(N__13135));
    LocalMux I__989 (
            .O(N__13135),
            .I(N__13132));
    Odrv4 I__988 (
            .O(N__13132),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__987 (
            .O(N__13129),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ));
    CascadeMux I__986 (
            .O(N__13126),
            .I(\this_vga_signals.g3_1_cascade_ ));
    CascadeMux I__985 (
            .O(N__13123),
            .I(\this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_ ));
    CascadeMux I__984 (
            .O(N__13120),
            .I(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ));
    CascadeMux I__983 (
            .O(N__13117),
            .I(\this_vga_signals.g1_1_cascade_ ));
    CascadeMux I__982 (
            .O(N__13114),
            .I(\this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_ ));
    defparam IN_MUX_bfv_24_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_24_21_0_));
    defparam IN_MUX_bfv_24_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_24_22_0_ (
            .carryinitin(un1_M_this_ext_address_q_cry_7),
            .carryinitout(bfn_24_22_0_));
    defparam IN_MUX_bfv_21_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_20_0_));
    defparam IN_MUX_bfv_21_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_21_0_ (
            .carryinitin(\this_ppu.un1_oam_data_1_cry_7 ),
            .carryinitout(bfn_21_21_0_));
    defparam IN_MUX_bfv_21_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_23_0_));
    defparam IN_MUX_bfv_21_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_24_0_ (
            .carryinitin(\this_ppu.un1_M_voffset_d_cry_7 ),
            .carryinitout(bfn_21_24_0_));
    defparam IN_MUX_bfv_20_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_24_0_));
    defparam IN_MUX_bfv_22_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_21_0_));
    defparam IN_MUX_bfv_22_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_22_0_ (
            .carryinitin(\this_ppu.un1_M_oam_cache_read_data_3_cry_7 ),
            .carryinitout(bfn_22_22_0_));
    defparam IN_MUX_bfv_20_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_19_0_));
    defparam IN_MUX_bfv_20_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_20_0_ (
            .carryinitin(\this_ppu.un1_M_oam_cache_read_data_2_cry_7 ),
            .carryinitout(bfn_20_20_0_));
    defparam IN_MUX_bfv_22_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_18_0_));
    defparam IN_MUX_bfv_22_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_19_0_ (
            .carryinitin(\this_ppu.un1_M_hoffset_q_cry_7 ),
            .carryinitout(bfn_22_19_0_));
    defparam IN_MUX_bfv_19_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_17_0_));
    defparam IN_MUX_bfv_19_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_18_0_ (
            .carryinitin(\this_ppu.un1_M_hoffset_d_cry_7 ),
            .carryinitout(bfn_19_18_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_3_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_9_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_21_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_22_0_));
    defparam IN_MUX_bfv_22_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_24_0_));
    defparam IN_MUX_bfv_22_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_25_0_ (
            .carryinitin(\this_ppu.un1_M_voffset_q_cry_7 ),
            .carryinitout(bfn_22_25_0_));
    defparam IN_MUX_bfv_21_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_18_0_));
    defparam IN_MUX_bfv_21_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_19_0_ (
            .carryinitin(\this_ppu.un1_M_hoffset_q_2_cry_7 ),
            .carryinitout(bfn_21_19_0_));
    defparam IN_MUX_bfv_21_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_17_0_));
    defparam IN_MUX_bfv_19_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_13_0_));
    defparam IN_MUX_bfv_19_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_14_0_ (
            .carryinitin(un1_M_this_spr_address_q_cry_7),
            .carryinitout(bfn_19_14_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_9_22_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNIR1G77_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__13264),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_935_0_g ));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNI67JU6_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__19210),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1212_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__23974),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__22600),
            .GLOBALBUFFEROUTPUT(N_504_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI93SL3_6_LC_1_8_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI93SL3_6_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI93SL3_6_LC_1_8_3 .LUT_INIT=16'b0011110001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI93SL3_6_LC_1_8_3  (
            .in0(N__17404),
            .in1(N__16133),
            .in2(N__13408),
            .in3(N__16603),
            .lcout(\this_vga_signals.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIDHDA1_1_LC_1_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIDHDA1_1_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIDHDA1_1_LC_1_9_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIDHDA1_1_LC_1_9_6  (
            .in0(N__15673),
            .in1(N__15400),
            .in2(_gnd_net_),
            .in3(N__15599),
            .lcout(\this_vga_signals.vaddress_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNI0SND1_LC_1_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNI0SND1_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_RNI0SND1_LC_1_9_7 .LUT_INIT=16'b0110111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_RNI0SND1_LC_1_9_7  (
            .in0(N__15205),
            .in1(N__16580),
            .in2(N__13597),
            .in3(N__13563),
            .lcout(\this_vga_signals.N_32_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_LC_1_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_LC_1_10_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_a5_1_LC_1_10_0  (
            .in0(N__15856),
            .in1(N__14695),
            .in2(N__16858),
            .in3(N__14582),
            .lcout(\this_vga_signals.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_1_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_1_10_1 .LUT_INIT=16'b1001011101101101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_1_10_1  (
            .in0(N__13709),
            .in1(N__16841),
            .in2(N__17576),
            .in3(N__14285),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_LC_1_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_LC_1_10_2 .LUT_INIT=16'b1110110110000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_LC_1_10_2  (
            .in0(N__14959),
            .in1(N__15490),
            .in2(N__13117),
            .in3(N__15620),
            .lcout(\this_vga_signals.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_1_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_1_10_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_a0_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__17475),
            .in2(_gnd_net_),
            .in3(N__16836),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_1_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_1_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_1_10_5  (
            .in0(N__17530),
            .in1(N__16840),
            .in2(_gnd_net_),
            .in3(N__14284),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_1_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_1_10_6 .LUT_INIT=16'b0010001000100011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_1_10_6  (
            .in0(N__14958),
            .in1(N__14075),
            .in2(N__13114),
            .in3(N__13710),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_1_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_2_LC_1_10_7 .LUT_INIT=16'b1111111101111011;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_2_LC_1_10_7  (
            .in0(N__13429),
            .in1(N__15480),
            .in2(N__13129),
            .in3(N__13853),
            .lcout(\this_vga_signals.g3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_1_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_10_LC_1_11_0 .LUT_INIT=16'b0111111010110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_10_LC_1_11_0  (
            .in0(N__16846),
            .in1(N__17390),
            .in2(N__17569),
            .in3(N__14692),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_1_LC_1_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_1_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_1_LC_1_11_1 .LUT_INIT=16'b0000000011101101;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_1_LC_1_11_1  (
            .in0(N__14282),
            .in1(N__17516),
            .in2(N__16859),
            .in3(N__13704),
            .lcout(),
            .ltout(\this_vga_signals.g3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_1_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_1_11_2 .LUT_INIT=16'b0011001011111010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_1_11_2  (
            .in0(N__14953),
            .in1(N__13138),
            .in2(N__13126),
            .in3(N__14283),
            .lcout(\this_vga_signals.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_rn_LC_1_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_rn_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_rn_LC_1_11_3 .LUT_INIT=16'b0000100110010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_rn_LC_1_11_3  (
            .in0(N__15765),
            .in1(N__15838),
            .in2(N__13795),
            .in3(N__14570),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_2_mb_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_mb_LC_1_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_mb_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_mb_LC_1_11_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_mb_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__14691),
            .in2(N__13123),
            .in3(N__13639),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_1_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14386),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40414),
            .ce(N__16293),
            .sr(N__16261));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_1_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_1_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_1_11_6  (
            .in0(N__17512),
            .in1(N__16842),
            .in2(_gnd_net_),
            .in3(N__14281),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axb1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_1_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_1_11_7 .LUT_INIT=16'b0011110010010011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_x4_LC_1_11_7  (
            .in0(N__17520),
            .in1(N__14952),
            .in2(N__13120),
            .in3(N__13703),
            .lcout(\this_vga_signals.if_N_9_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_i_o2_LC_1_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_i_o2_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_i_o2_LC_1_12_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_i_o2_LC_1_12_0  (
            .in0(N__14265),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16778),
            .lcout(\this_vga_signals.g2_1_0 ),
            .ltout(\this_vga_signals.g2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_1_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_LC_1_12_1 .LUT_INIT=16'b1010101011101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_LC_1_12_1  (
            .in0(N__14950),
            .in1(N__17590),
            .in2(N__13159),
            .in3(N__13708),
            .lcout(),
            .ltout(\this_vga_signals.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_1_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_1_12_2 .LUT_INIT=16'b0110010110011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_a2_LC_1_12_2  (
            .in0(N__13653),
            .in1(N__14065),
            .in2(N__13156),
            .in3(N__13986),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_1_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_1_12_3 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_1_LC_1_12_3  (
            .in0(N__15837),
            .in1(N__15772),
            .in2(_gnd_net_),
            .in3(N__14264),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_ac0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_1_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_12_LC_1_12_4 .LUT_INIT=16'b0000000011001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_12_LC_1_12_4  (
            .in0(N__13706),
            .in1(N__14951),
            .in2(N__13153),
            .in3(N__14064),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_1_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_0_LC_1_12_5 .LUT_INIT=16'b0011001000110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_0_LC_1_12_5  (
            .in0(N__16779),
            .in1(N__13705),
            .in2(N__17598),
            .in3(N__14266),
            .lcout(\this_vga_signals.g3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_0_LC_1_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_0_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_0_LC_1_12_6 .LUT_INIT=16'b0111111111101111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_0_LC_1_12_6  (
            .in0(N__17389),
            .in1(N__14696),
            .in2(N__13150),
            .in3(N__14583),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_1_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_1_12_7 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_1_12_7  (
            .in0(N__14063),
            .in1(N__13707),
            .in2(N__14973),
            .in3(N__13746),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_LC_1_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_LC_1_13_0 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_LC_1_13_0  (
            .in0(N__17392),
            .in1(N__17563),
            .in2(N__16822),
            .in3(N__14705),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_1_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_1_13_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14302),
            .in3(N__16774),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_1_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_LC_1_13_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_LC_1_13_2  (
            .in0(N__13970),
            .in1(_gnd_net_),
            .in2(N__13183),
            .in3(N__15627),
            .lcout(\this_vga_signals.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_0_LC_1_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_0_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_0_LC_1_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_0_LC_1_13_3  (
            .in0(N__17564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13969),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(\this_vga_signals.g1_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_x0_LC_1_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_x0_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_x0_LC_1_13_4 .LUT_INIT=16'b1111101111110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_x0_LC_1_13_4  (
            .in0(N__13971),
            .in1(N__15476),
            .in2(N__13180),
            .in3(N__14011),
            .lcout(\this_vga_signals.g3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_1_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_1_13_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_1_13_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__14356),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40428),
            .ce(N__16292),
            .sr(N__16263));
    defparam \this_vga_signals.un5_vaddress_g3_x1_LC_1_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_x1_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_x1_LC_1_13_6 .LUT_INIT=16'b0110111111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_x1_LC_1_13_6  (
            .in0(N__13972),
            .in1(N__14012),
            .in2(N__15520),
            .in3(N__13177),
            .lcout(\this_vga_signals.g3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_1_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_1_13_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__14355),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40428),
            .ce(N__16292),
            .sr(N__16263));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_1_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_1_14_0 .LUT_INIT=16'b0001011101001101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_c2_LC_1_14_0  (
            .in0(N__17567),
            .in1(N__13887),
            .in2(N__15513),
            .in3(N__13976),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1NB793_6_LC_1_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1NB793_6_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI1NB793_6_LC_1_14_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI1NB793_6_LC_1_14_1  (
            .in0(N__13171),
            .in1(N__14118),
            .in2(N__13162),
            .in3(N__13278),
            .lcout(\this_vga_signals.g2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_1_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_1_14_2 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_1_LC_1_14_2  (
            .in0(N__17566),
            .in1(N__13886),
            .in2(N__15512),
            .in3(N__13974),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_LC_1_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_LC_1_14_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_LC_1_14_3  (
            .in0(N__13852),
            .in1(N__13327),
            .in2(N__14748),
            .in3(N__13195),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axb1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_1_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_1_14_4 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_1_14_4  (
            .in0(N__15688),
            .in1(N__13258),
            .in2(N__13249),
            .in3(N__13801),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBN8KM1_4_LC_1_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBN8KM1_4_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBN8KM1_4_LC_1_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBN8KM1_4_LC_1_14_5  (
            .in0(N__13975),
            .in1(N__13246),
            .in2(N__13898),
            .in3(N__17568),
            .lcout(\this_vga_signals.vaddress_m2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_1_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m1_0_LC_1_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m1_0_LC_1_14_6  (
            .in0(N__17565),
            .in1(N__13973),
            .in2(_gnd_net_),
            .in3(N__13885),
            .lcout(\this_vga_signals.if_m1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_1_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_1_15_0 .LUT_INIT=16'b1011001000001111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m8_0_m2_LC_1_15_0  (
            .in0(N__15632),
            .in1(N__13234),
            .in2(N__15516),
            .in3(N__13225),
            .lcout(\this_vga_signals.mult1_un68_sum_c3 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_1_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_3_LC_1_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_3_LC_1_15_1  (
            .in0(N__15008),
            .in1(N__13912),
            .in2(N__13219),
            .in3(N__13194),
            .lcout(\this_vga_signals.g2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_1_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_LC_1_15_2 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_LC_1_15_2  (
            .in0(N__13216),
            .in1(N__14125),
            .in2(N__15517),
            .in3(N__14020),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_1_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_1_15_3 .LUT_INIT=16'b1000010000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_1_15_3  (
            .in0(N__13207),
            .in1(N__15687),
            .in2(N__13201),
            .in3(N__14189),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_1_LC_1_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_1_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_1_LC_1_15_4 .LUT_INIT=16'b0011001101101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_1_LC_1_15_4  (
            .in0(N__17585),
            .in1(N__15621),
            .in2(N__15515),
            .in3(N__13990),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axb1_3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_LC_1_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_LC_1_15_5 .LUT_INIT=16'b0001111001111000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb1_3_1_LC_1_15_5  (
            .in0(N__15505),
            .in1(N__17586),
            .in2(N__13198),
            .in3(N__13900),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_1_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_1_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_LC_1_15_6  (
            .in0(N__13899),
            .in1(N__15007),
            .in2(N__14980),
            .in3(N__13991),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_1_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_14_LC_1_15_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_14_LC_1_15_7  (
            .in0(N__13992),
            .in1(N__15498),
            .in2(N__13369),
            .in3(N__15633),
            .lcout(\this_vga_signals.g0_0_0_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_1_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_4_LC_1_16_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_4_LC_1_16_0  (
            .in0(N__13612),
            .in1(N__14223),
            .in2(N__13357),
            .in3(N__13325),
            .lcout(),
            .ltout(\this_vga_signals.g1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_1_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_1_16_1 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_1_16_1  (
            .in0(N__15052),
            .in1(N__14744),
            .in2(N__13345),
            .in3(N__14169),
            .lcout(\this_vga_signals.if_i4_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_1_16_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_1_16_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_1_16_2  (
            .in0(N__16915),
            .in1(N__17002),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNILB7N84_2_LC_1_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNILB7N84_2_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNILB7N84_2_LC_1_16_3 .LUT_INIT=16'b0001010011101011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNILB7N84_2_LC_1_16_3  (
            .in0(N__13326),
            .in1(N__15637),
            .in2(N__15519),
            .in3(N__13312),
            .lcout(\this_vga_signals.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_1_16_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_1_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13303),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40449),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_1_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_1_16_6 .LUT_INIT=16'b1000110101001110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_1_16_6  (
            .in0(N__14098),
            .in1(N__13291),
            .in2(N__15518),
            .in3(N__13282),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIR1G77_9_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(N__20064),
            .in2(_gnd_net_),
            .in3(N__16267),
            .lcout(\this_vga_signals.N_935_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.port_data_rw_0_i_LC_1_18_1 .C_ON=1'b0;
    defparam \this_ppu.port_data_rw_0_i_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.port_data_rw_0_i_LC_1_18_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_ppu.port_data_rw_0_i_LC_1_18_1  (
            .in0(N__29223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32217),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQPR1_7_LC_2_8_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQPR1_7_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIUQPR1_7_LC_2_8_3 .LUT_INIT=16'b1011010001001011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIUQPR1_7_LC_2_8_3  (
            .in0(N__17570),
            .in1(N__16860),
            .in2(N__14134),
            .in3(N__16708),
            .lcout(\this_vga_signals.g2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_2_8_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_2_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__16976),
            .in2(_gnd_net_),
            .in3(N__17059),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_2_8_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_2_8_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_2_8_6  (
            .in0(N__17020),
            .in1(_gnd_net_),
            .in2(N__16992),
            .in3(_gnd_net_),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_0_9_LC_2_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_0_9_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_0_9_LC_2_9_0 .LUT_INIT=16'b0001101000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_0_9_LC_2_9_0  (
            .in0(N__13447),
            .in1(N__14415),
            .in2(N__13468),
            .in3(N__15139),
            .lcout(\this_vga_signals.SUM_2_i_i_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_2_9_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_2_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_2_9_1  (
            .in0(N__15918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_2_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_2_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_2_9_2  (
            .in0(N__16313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_2_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15869),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_N_2L1_LC_2_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_N_2L1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_N_2L1_LC_2_9_4 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_N_2L1_LC_2_9_4  (
            .in0(N__14430),
            .in1(N__13506),
            .in2(N__13542),
            .in3(N__14414),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_2_2_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_2_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14375),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_2_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_2_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14452),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_2_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_2_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14346),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40385),
            .ce(N__16298),
            .sr(N__16255));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_9_LC_2_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_9_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_9_LC_2_10_0 .LUT_INIT=16'b1010011110101111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIRK3H_9_LC_2_10_0  (
            .in0(N__15136),
            .in1(N__13445),
            .in2(N__13467),
            .in3(N__14413),
            .lcout(\this_vga_signals.SUM_2_i_i_1_0_3 ),
            .ltout(\this_vga_signals.SUM_2_i_i_1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x0_LC_2_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x0_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x0_LC_2_10_1 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x0_LC_2_10_1  (
            .in0(N__15184),
            .in1(N__15255),
            .in2(N__13450),
            .in3(N__16565),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_2_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_2_10_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_0_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13541),
            .in3(N__13504),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_x1_LC_2_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_x1_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_x1_LC_2_10_3 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_x1_LC_2_10_3  (
            .in0(N__13446),
            .in1(N__15256),
            .in2(N__15314),
            .in3(N__15137),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_2_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_ns_LC_2_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_ns_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_ns_LC_2_10_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_ns_LC_2_10_4  (
            .in0(N__16566),
            .in1(_gnd_net_),
            .in2(N__13432),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_2_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_2_LC_2_10_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_2_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13993),
            .in3(N__17529),
            .lcout(\this_vga_signals.g1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x1_LC_2_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x1_LC_2_10_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x1_LC_2_10_6  (
            .in0(N__15138),
            .in1(N__13505),
            .in2(N__15270),
            .in3(N__15305),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_ns_LC_2_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_ns_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_ns_LC_2_10_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_ns_LC_2_10_7  (
            .in0(N__13570),
            .in1(_gnd_net_),
            .in2(N__13600),
            .in3(N__13534),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_ns ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_ns_LC_2_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_ns_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_ns_LC_2_11_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_ns_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__13596),
            .in2(N__13579),
            .in3(N__13549),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x0_LC_2_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x0_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x0_LC_2_11_1 .LUT_INIT=16'b0000010000000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a3_x0_LC_2_11_1  (
            .in0(N__15253),
            .in1(N__15140),
            .in2(N__15313),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_2_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_2_11_2 .LUT_INIT=16'b0110000110010100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb2_LC_2_11_2  (
            .in0(N__14569),
            .in1(N__13794),
            .in2(N__13633),
            .in3(N__14693),
            .lcout(\this_vga_signals.mult1_un54_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x1_LC_2_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x1_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x1_LC_2_11_3 .LUT_INIT=16'b1111101000111001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_axb1_x1_LC_2_11_3  (
            .in0(N__15183),
            .in1(N__15260),
            .in2(N__13564),
            .in3(N__16567),
            .lcout(\this_vga_signals.mult1_un40_sum_axb1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_x1_LC_2_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_x1_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_x1_LC_2_11_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_x1_LC_2_11_4  (
            .in0(N__15141),
            .in1(N__13543),
            .in2(N__15200),
            .in3(N__15254),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_ns_LC_2_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_ns_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_ns_LC_2_11_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_0_a0_ns_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13513),
            .in3(N__13510),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_0_a0_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_2_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_2_11_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_2_11_6  (
            .in0(N__13486),
            .in1(N__14458),
            .in2(N__13480),
            .in3(N__13477),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_2_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_2_11_7 .LUT_INIT=16'b1000101101010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_ac0_3_LC_2_11_7  (
            .in0(N__13793),
            .in1(N__13628),
            .in2(N__13471),
            .in3(N__14568),
            .lcout(\this_vga_signals.mult1_un47_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_sn_LC_2_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_sn_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_sn_LC_2_12_0 .LUT_INIT=16'b0010000100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_2_mb_sn_LC_2_12_0  (
            .in0(N__15763),
            .in1(N__13632),
            .in2(N__15839),
            .in3(N__14565),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_2_mb_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_2_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_2_12_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_2_12_1  (
            .in0(N__15821),
            .in1(N__15757),
            .in2(_gnd_net_),
            .in3(N__15263),
            .lcout(\this_vga_signals.r_N_4_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_2_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_2_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_2_12_2  (
            .in0(N__14382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40419),
            .ce(N__16294),
            .sr(N__16262));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_2_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_2_12_3 .LUT_INIT=16'b1000100001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_2_12_3  (
            .in0(N__15823),
            .in1(N__15761),
            .in2(_gnd_net_),
            .in3(N__15261),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_2_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_2_12_4 .LUT_INIT=16'b0101010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_0_LC_2_12_4  (
            .in0(N__15262),
            .in1(_gnd_net_),
            .in2(N__15773),
            .in3(N__15822),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1_0 ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_2_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_2_12_5 .LUT_INIT=16'b0010000000010100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_4_LC_2_12_5  (
            .in0(N__14566),
            .in1(N__14694),
            .in2(N__13615),
            .in3(N__13792),
            .lcout(\this_vga_signals.mult1_un54_sum_ac0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_0_LC_2_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_0_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_0_LC_2_12_6 .LUT_INIT=16'b0111111010011111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_1_0_LC_2_12_6  (
            .in0(N__15762),
            .in1(N__15824),
            .in2(N__17403),
            .in3(N__14690),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_3_LC_2_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_3_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_3_LC_2_12_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_a5_1_3_LC_2_12_7  (
            .in0(N__14567),
            .in1(N__17399),
            .in2(_gnd_net_),
            .in3(N__15764),
            .lcout(\this_vga_signals.g0_0_i_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_2_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_2_13_0 .LUT_INIT=16'b0000000011001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_2_13_0  (
            .in0(N__13747),
            .in1(N__14974),
            .in2(N__13717),
            .in3(N__14062),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_2_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_2_13_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_3_LC_2_13_1  (
            .in0(N__13968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17572),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_3_LC_2_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_3_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_3_LC_2_13_2 .LUT_INIT=16'b1111111101111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_3_LC_2_13_2  (
            .in0(N__15491),
            .in1(N__13813),
            .in2(N__13807),
            .in3(N__13851),
            .lcout(\this_vga_signals.g3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_2_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_2_13_3 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_2_13_3  (
            .in0(N__14061),
            .in1(N__14960),
            .in2(N__13748),
            .in3(N__13711),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_2_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_2_13_4 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb2_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__14013),
            .in2(N__13804),
            .in3(N__13967),
            .lcout(\this_vga_signals.mult1_un61_sum_axb2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_0_LC_2_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_0_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_0_LC_2_13_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_0_LC_2_13_5  (
            .in0(N__16046),
            .in1(N__14485),
            .in2(_gnd_net_),
            .in3(N__14813),
            .lcout(\this_vga_signals.g0_0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_2_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_2_13_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_LC_2_13_6  (
            .in0(N__14592),
            .in1(N__13791),
            .in2(N__14301),
            .in3(N__13762),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_2_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_2_13_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_1_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13753),
            .in3(N__17571),
            .lcout(\this_vga_signals.g1_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_1_LC_2_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_1_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_1_LC_2_14_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axbxc3_1_1_LC_2_14_0  (
            .in0(N__13715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13749),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_2_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_2_14_1 .LUT_INIT=16'b0000110000001101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_2_14_1  (
            .in0(N__13750),
            .in1(N__14961),
            .in2(N__14082),
            .in3(N__13716),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_0_LC_2_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_0_LC_2_14_2 .LUT_INIT=16'b1100110010000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_0_LC_2_14_2  (
            .in0(N__13985),
            .in1(N__14626),
            .in2(N__13660),
            .in3(N__13657),
            .lcout(\this_vga_signals.g0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_6_LC_2_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_6_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_6_LC_2_14_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_6_LC_2_14_3  (
            .in0(N__14293),
            .in1(N__14119),
            .in2(N__16531),
            .in3(N__16161),
            .lcout(\this_vga_signals.g0_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_2_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_2_14_4 .LUT_INIT=16'b1010010110100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_2_14_4  (
            .in0(N__14089),
            .in1(N__14969),
            .in2(N__14083),
            .in3(N__14032),
            .lcout(\this_vga_signals.N_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_4_LC_2_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_4_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_4_LC_2_14_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_4_LC_2_14_5  (
            .in0(N__14014),
            .in1(N__13891),
            .in2(_gnd_net_),
            .in3(N__13984),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_0_0_LC_2_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_0_0_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_0_0_LC_2_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_0_0_LC_2_14_6  (
            .in0(N__14962),
            .in1(N__16780),
            .in2(_gnd_net_),
            .in3(N__14292),
            .lcout(\this_vga_signals.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_ns_LC_2_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_ns_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_ns_LC_2_14_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_ns_LC_2_14_7  (
            .in0(N__13906),
            .in1(N__13892),
            .in2(_gnd_net_),
            .in3(N__13861),
            .lcout(\this_vga_signals.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_LC_2_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_LC_2_15_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_LC_2_15_0  (
            .in0(N__13855),
            .in1(N__14217),
            .in2(N__15040),
            .in3(N__14738),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_2_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_2_15_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_2_15_1  (
            .in0(N__14979),
            .in1(N__15013),
            .in2(N__16855),
            .in3(N__14304),
            .lcout(\this_vga_signals.g0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_2_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_2_15_2 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_LC_2_15_2  (
            .in0(N__13854),
            .in1(N__14599),
            .in2(N__13822),
            .in3(N__14812),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_2_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_2_15_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_2_15_3  (
            .in0(N__14740),
            .in1(N__14227),
            .in2(N__14323),
            .in3(N__14320),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI7RTI411_2_LC_2_15_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI7RTI411_2_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI7RTI411_2_LC_2_15_4 .LUT_INIT=16'b0101010110011010;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI7RTI411_2_LC_2_15_4  (
            .in0(N__14191),
            .in1(N__15610),
            .in2(N__14314),
            .in3(N__14311),
            .lcout(\this_vga_signals.vaddress_m6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_0_a2_3_LC_2_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_a2_3_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_a2_3_LC_2_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_0_a2_3_LC_2_15_5  (
            .in0(N__14218),
            .in1(N__16823),
            .in2(_gnd_net_),
            .in3(N__14303),
            .lcout(\this_vga_signals.g0_6_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_0_a2_2_LC_2_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_0_a2_2_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_0_a2_2_LC_2_15_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_0_a2_2_LC_2_15_6  (
            .in0(N__14305),
            .in1(N__14219),
            .in2(N__16854),
            .in3(N__14739),
            .lcout(),
            .ltout(\this_vga_signals.g3_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_2_15_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_2_15_7 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_2_15_7  (
            .in0(N__15609),
            .in1(N__14614),
            .in2(N__14194),
            .in3(N__14190),
            .lcout(\this_vga_signals.mult1_un75_sum_ac0_3_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_2_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_2_16_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_9_LC_2_16_1  (
            .in0(N__20510),
            .in1(N__17595),
            .in2(N__16856),
            .in3(N__16408),
            .lcout(\this_vga_signals.vsync_1_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIGAFCKA_2_LC_2_16_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIGAFCKA_2_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIGAFCKA_2_LC_2_16_3 .LUT_INIT=16'b1001110011000110;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIGAFCKA_2_LC_2_16_3  (
            .in0(N__15631),
            .in1(N__14176),
            .in2(N__15514),
            .in3(N__14170),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_N_3_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI0FQEQV_2_LC_2_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI0FQEQV_2_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI0FQEQV_2_LC_2_16_4 .LUT_INIT=16'b1000101101000111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI0FQEQV_2_LC_2_16_4  (
            .in0(N__14158),
            .in1(N__14152),
            .in2(N__14146),
            .in3(N__14143),
            .lcout(\this_vga_signals.M_vcounter_q_RNI0FQEQVZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_6_LC_3_8_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_6_LC_3_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICSHP_6_LC_3_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICSHP_6_LC_3_8_5  (
            .in0(_gnd_net_),
            .in1(N__15380),
            .in2(_gnd_net_),
            .in3(N__17393),
            .lcout(\this_vga_signals.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_3_9_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_3_9_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_3_9_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_3_9_0  (
            .in0(N__20068),
            .in1(N__15339),
            .in2(N__19894),
            .in3(N__19890),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_3_9_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__40378),
            .ce(),
            .sr(N__16254));
    defparam \this_vga_signals.M_vcounter_q_1_LC_3_9_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_3_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_3_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_3_9_1  (
            .in0(N__20070),
            .in1(N__15672),
            .in2(_gnd_net_),
            .in3(N__14395),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__40378),
            .ce(),
            .sr(N__16254));
    defparam \this_vga_signals.M_vcounter_q_2_LC_3_9_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_3_9_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_3_9_2  (
            .in0(N__20069),
            .in1(N__15576),
            .in2(_gnd_net_),
            .in3(N__14392),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__40378),
            .ce(),
            .sr(N__16254));
    defparam \this_vga_signals.M_vcounter_q_3_LC_3_9_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_3_9_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_3_9_3  (
            .in0(N__20071),
            .in1(N__15422),
            .in2(_gnd_net_),
            .in3(N__14389),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__40378),
            .ce(),
            .sr(N__16254));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_3_9_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_3_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_3_9_4  (
            .in0(_gnd_net_),
            .in1(N__17596),
            .in2(_gnd_net_),
            .in3(N__14359),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_3_9_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_3_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_3_9_5  (
            .in0(_gnd_net_),
            .in1(N__16857),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_3_9_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_3_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_3_9_6  (
            .in0(_gnd_net_),
            .in1(N__17394),
            .in2(_gnd_net_),
            .in3(N__14332),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_3_9_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_3_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_3_9_7  (
            .in0(_gnd_net_),
            .in1(N__16706),
            .in2(_gnd_net_),
            .in3(N__14329),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_3_10_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_3_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(_gnd_net_),
            .in3(N__14326),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_3_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_3_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__20484),
            .in2(_gnd_net_),
            .in3(N__14473),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_3_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_3_10_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_3_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_9_rep1_esr_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15917),
            .lcout(\this_vga_signals.M_vcounter_q_9_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40386),
            .ce(N__16299),
            .sr(N__16256));
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_3_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_3_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_8_rep1_esr_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14450),
            .lcout(\this_vga_signals.M_vcounter_q_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40386),
            .ce(N__16299),
            .sr(N__16256));
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_3_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_3_LC_3_11_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_3_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__14954),
            .in2(_gnd_net_),
            .in3(N__15012),
            .lcout(\this_vga_signals.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_LC_3_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_LC_3_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_LC_3_11_3 .LUT_INIT=16'b1000101111001101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_2_2_LC_3_11_3  (
            .in0(N__16376),
            .in1(N__15185),
            .in2(N__14470),
            .in3(N__15306),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_3_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_3_11_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_3_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_7_rep1_esr_LC_3_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16320),
            .lcout(\this_vga_signals.M_vcounter_q_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40398),
            .ce(N__16296),
            .sr(N__16258));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_3_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_3_11_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_3_11_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_3_11_5  (
            .in0(_gnd_net_),
            .in1(N__14451),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_vga_signals_M_vcounter_q_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40398),
            .ce(N__16296),
            .sr(N__16258));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_3_11_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_3_11_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_3_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_3_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15876),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40398),
            .ce(N__16296),
            .sr(N__16258));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_1_a0_1_LC_3_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_1_a0_1_LC_3_12_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_1_a0_1_LC_3_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_1_a0_1_LC_3_12_0  (
            .in0(_gnd_net_),
            .in1(N__14434),
            .in2(_gnd_net_),
            .in3(N__14419),
            .lcout(),
            .ltout(\this_vga_signals.N_1_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_1_LC_3_12_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_1_LC_3_12_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_1_LC_3_12_1 .LUT_INIT=16'b0110011111101111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_1_LC_3_12_1  (
            .in0(N__15316),
            .in1(N__16688),
            .in2(N__14512),
            .in3(N__15699),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_c2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_3_12_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_3_12_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_3_12_2 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_LC_3_12_2  (
            .in0(N__16594),
            .in1(N__14479),
            .in2(N__14509),
            .in3(N__14500),
            .lcout(\this_vga_signals.mult1_un40_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un40_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_3_12_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_3_12_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_3_12_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_3_12_3  (
            .in0(N__15934),
            .in1(_gnd_net_),
            .in2(N__14506),
            .in3(N__16156),
            .lcout(\this_vga_signals.N_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIOKSG_LC_3_12_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIOKSG_LC_3_12_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIOKSG_LC_3_12_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIOKSG_LC_3_12_4  (
            .in0(_gnd_net_),
            .in1(N__16378),
            .in2(_gnd_net_),
            .in3(N__15268),
            .lcout(\this_vga_signals.vaddress_m2_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_3_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_3_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_3_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_3_12_5  (
            .in0(N__16179),
            .in1(N__16155),
            .in2(_gnd_net_),
            .in3(N__16097),
            .lcout(\this_vga_signals.g0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_1_0_LC_3_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_1_0_LC_3_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_1_0_LC_3_12_6 .LUT_INIT=16'b0110011011011101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_1_0_LC_3_12_6  (
            .in0(N__15198),
            .in1(N__16377),
            .in2(_gnd_net_),
            .in3(N__15315),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_c2_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_LC_3_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_LC_3_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_LC_3_12_7 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_c2_2_LC_3_12_7  (
            .in0(N__15269),
            .in1(_gnd_net_),
            .in2(N__14503),
            .in3(N__16593),
            .lcout(\this_vga_signals.mult1_un40_sum_c2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_3_13_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_3_13_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_3_13_0 .LUT_INIT=16'b0100010111101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_5_LC_3_13_0  (
            .in0(N__14494),
            .in1(N__14591),
            .in2(N__17251),
            .in3(N__16024),
            .lcout(\this_vga_signals.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_LC_3_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_LC_3_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_LC_3_13_1 .LUT_INIT=16'b0111000001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_LC_3_13_1  (
            .in0(N__15201),
            .in1(N__16590),
            .in2(N__15109),
            .in3(N__15271),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_3_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_3_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_3_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a0_2_LC_3_13_2  (
            .in0(N__16591),
            .in1(N__14590),
            .in2(N__17380),
            .in3(N__14706),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_LC_3_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_LC_3_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_LC_3_13_3 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_a5_LC_3_13_3  (
            .in0(N__14707),
            .in1(N__14647),
            .in2(N__16853),
            .in3(N__15888),
            .lcout(),
            .ltout(\this_vga_signals.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_3_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_3_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_3_13_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_2_LC_3_13_4  (
            .in0(N__15889),
            .in1(N__14641),
            .in2(N__14629),
            .in3(N__16023),
            .lcout(\this_vga_signals.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_8_LC_3_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_8_LC_3_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_8_LC_3_13_5 .LUT_INIT=16'b0101111101111110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_8_LC_3_13_5  (
            .in0(N__16705),
            .in1(N__16592),
            .in2(N__16407),
            .in3(N__17350),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_3_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_3_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_3_13_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_0_LC_3_13_7  (
            .in0(N__16180),
            .in1(N__16160),
            .in2(_gnd_net_),
            .in3(N__16099),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_3_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_1_0_LC_3_14_0 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_1_0_LC_3_14_0  (
            .in0(N__14814),
            .in1(N__14878),
            .in2(N__16003),
            .in3(N__14620),
            .lcout(\this_vga_signals.g3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_3_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_3_14_1 .LUT_INIT=16'b0010000000101010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_0_2_LC_3_14_1  (
            .in0(N__16056),
            .in1(N__16071),
            .in2(N__14608),
            .in3(N__16026),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_1_LC_3_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_1_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_1_LC_3_14_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_1_LC_3_14_2  (
            .in0(N__17594),
            .in1(N__17345),
            .in2(_gnd_net_),
            .in3(N__14593),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_3_14_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_3_14_3 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_3_14_3  (
            .in0(N__16055),
            .in1(N__14524),
            .in2(N__14515),
            .in3(N__16025),
            .lcout(\this_vga_signals.g0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_0_LC_3_14_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_0_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_0_LC_3_14_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un75_sum_axb2_0_LC_3_14_4  (
            .in0(N__15423),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15597),
            .lcout(\this_vga_signals.mult1_un75_sum_axb2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_14_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_14_5  (
            .in0(_gnd_net_),
            .in1(N__17113),
            .in2(_gnd_net_),
            .in3(N__16993),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_7_LC_3_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_7_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI87V41_7_LC_3_14_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI87V41_7_LC_3_14_6  (
            .in0(N__16707),
            .in1(N__17346),
            .in2(_gnd_net_),
            .in3(N__15598),
            .lcout(\this_vga_signals.vsync_1_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g3_0_1_LC_3_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g3_0_1_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g3_0_1_LC_3_14_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g3_0_1_LC_3_14_7  (
            .in0(_gnd_net_),
            .in1(N__15006),
            .in2(_gnd_net_),
            .in3(N__14978),
            .lcout(\this_vga_signals.g3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_3_15_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_9_LC_3_15_0 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_9_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__14713),
            .in2(N__14872),
            .in3(N__14863),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_c3_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIU4E93J3_8_LC_3_15_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIU4E93J3_8_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIU4E93J3_8_LC_3_15_1 .LUT_INIT=16'b0010100010000010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIU4E93J3_8_LC_3_15_1  (
            .in0(N__15988),
            .in1(N__14854),
            .in2(N__14848),
            .in3(N__14845),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_3_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_13_LC_3_15_2 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_13_LC_3_15_2  (
            .in0(N__14815),
            .in1(N__14791),
            .in2(N__14782),
            .in3(N__14773),
            .lcout(),
            .ltout(\this_vga_signals.N_12_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_3_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_3_15_3 .LUT_INIT=16'b1110011110111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_3_15_3  (
            .in0(N__14767),
            .in1(N__14758),
            .in2(N__14752),
            .in3(N__14749),
            .lcout(\this_vga_signals.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_3_16_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_3_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_3_16_0  (
            .in0(N__17620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17001),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_3_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_3_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_3_16_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOLTE3_1_LC_3_16_5  (
            .in0(N__15680),
            .in1(N__15082),
            .in2(N__15073),
            .in3(N__15424),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_3_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_8_LC_3_16_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_8_LC_3_16_6  (
            .in0(_gnd_net_),
            .in1(N__15679),
            .in2(_gnd_net_),
            .in3(N__15340),
            .lcout(\this_vga_signals.if_N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_1_LC_4_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_4_8_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_4_8_6  (
            .in0(N__20077),
            .in1(N__18324),
            .in2(_gnd_net_),
            .in3(N__18376),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40353),
            .ce(),
            .sr(N__16515));
    defparam \this_vga_signals.M_hcounter_q_0_LC_4_8_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_4_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_4_8_7  (
            .in0(N__18325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20076),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40353),
            .ce(),
            .sr(N__16515));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_4_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_4_9_0 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_4_9_0  (
            .in0(N__18987),
            .in1(N__18185),
            .in2(_gnd_net_),
            .in3(N__18112),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_4_9_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_4_9_2 .LUT_INIT=16'b1100100000010011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axb1_LC_4_9_2  (
            .in0(N__18990),
            .in1(N__18187),
            .in2(N__18260),
            .in3(N__18234),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_4_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_4_9_3 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_4_9_3  (
            .in0(N__18815),
            .in1(N__19055),
            .in2(N__18918),
            .in3(N__18986),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_4_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_4_9_4 .LUT_INIT=16'b0010000011100000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_3_LC_4_9_4  (
            .in0(N__18988),
            .in1(N__18186),
            .in2(N__15043),
            .in3(N__18113),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_4_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_4_9_6 .LUT_INIT=16'b0101000001011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_1_LC_4_9_6  (
            .in0(N__18989),
            .in1(N__18114),
            .in2(N__18204),
            .in3(N__18233),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_4_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_4_9_7 .LUT_INIT=16'b0000000011010001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_4_9_7  (
            .in0(N__15721),
            .in1(N__18251),
            .in2(N__15715),
            .in3(N__15712),
            .lcout(\this_vga_signals.mult1_un61_sum_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_4_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_4_10_0 .LUT_INIT=16'b1001010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_4_10_0  (
            .in0(N__18809),
            .in1(N__19054),
            .in2(N__18917),
            .in3(N__18991),
            .lcout(\this_vga_signals.SUM_3_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_8_LC_4_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_8_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_8_LC_4_10_1 .LUT_INIT=16'b0010001001111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_0_8_LC_4_10_1  (
            .in0(N__16702),
            .in1(N__16380),
            .in2(N__17395),
            .in3(N__16601),
            .lcout(),
            .ltout(\this_vga_signals.vvisibility_i_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_9_LC_4_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_9_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_9_LC_4_10_2 .LUT_INIT=16'b0100000101010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_9_LC_4_10_2  (
            .in0(N__20483),
            .in1(N__16703),
            .in2(N__15706),
            .in3(N__15703),
            .lcout(N_825_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_4_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_4_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_8_LC_4_10_3  (
            .in0(N__17375),
            .in1(N__16698),
            .in2(N__16870),
            .in3(N__16379),
            .lcout(\this_vga_signals.M_lcounter_q_3_i_o2_2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_4_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_4_10_6 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_4_10_6  (
            .in0(N__15660),
            .in1(N__15550),
            .in2(N__15399),
            .in3(N__15335),
            .lcout(\this_vga_signals.N_822_0 ),
            .ltout(\this_vga_signals.N_822_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_4_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_4_10_7 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIBTPQ2_6_LC_4_10_7  (
            .in0(N__16869),
            .in1(N__17379),
            .in2(N__15319),
            .in3(N__17583),
            .lcout(this_vga_signals_un4_lvisibility_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_0_LC_4_11_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_0_LC_4_11_0 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_0_0_LC_4_11_0  (
            .in0(N__15307),
            .in1(N__15264),
            .in2(N__15199),
            .in3(N__15142),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_4_11_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_4_11_3 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_4_11_3  (
            .in0(N__17368),
            .in1(N__15844),
            .in2(_gnd_net_),
            .in3(N__15784),
            .lcout(),
            .ltout(\this_vga_signals.r_N_4_mux_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_1_9_LC_4_11_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_1_9_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_1_9_LC_4_11_4 .LUT_INIT=16'b1000011011110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI767P1_1_9_LC_4_11_4  (
            .in0(N__20443),
            .in1(N__16680),
            .in2(N__15937),
            .in3(N__16381),
            .lcout(\this_vga_signals.N_24_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_4_11_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_4_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI2UC41_0_LC_4_11_5  (
            .in0(N__18393),
            .in1(N__18535),
            .in2(N__18655),
            .in3(N__18331),
            .lcout(),
            .ltout(\this_vga_signals.un2_hsynclt6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_4_11_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_4_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIEVMV1_5_LC_4_11_6  (
            .in0(N__18142),
            .in1(N__18210),
            .in2(N__15925),
            .in3(N__19013),
            .lcout(\this_vga_signals.un2_hsynclt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_4_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_4_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15922),
            .lcout(this_vga_signals_M_vcounter_q_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40399),
            .ce(N__16297),
            .sr(N__16259));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI539J1_9_LC_4_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI539J1_9_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI539J1_9_LC_4_12_6 .LUT_INIT=16'b1001001011011101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI539J1_9_LC_4_12_6  (
            .in0(N__16686),
            .in1(N__15901),
            .in2(N__20479),
            .in3(N__16387),
            .lcout(),
            .ltout(\this_vga_signals.N_24_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_4_12_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_4_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_27_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__16154),
            .in2(N__15892),
            .in3(N__16096),
            .lcout(\this_vga_signals.N_4_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_4_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_4_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15880),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40408),
            .ce(N__16295),
            .sr(N__16260));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_0_LC_4_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_0_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a5_1_0_LC_4_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_a5_1_0_LC_4_13_2  (
            .in0(N__15783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17325),
            .lcout(\this_vga_signals.g0_0_i_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_4_13_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_4_13_3 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIDVUM_LC_4_13_3  (
            .in0(N__17326),
            .in1(N__15840),
            .in2(_gnd_net_),
            .in3(N__15782),
            .lcout(\this_vga_signals.r_N_4_mux ),
            .ltout(\this_vga_signals.r_N_4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_9_LC_4_13_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_9_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_9_LC_4_13_4 .LUT_INIT=16'b1000011011110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI767P1_9_LC_4_13_4  (
            .in0(N__20473),
            .in1(N__16682),
            .in2(N__16183),
            .in3(N__16398),
            .lcout(\this_vga_signals.N_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_0_9_LC_4_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_0_9_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI767P1_0_9_LC_4_13_5 .LUT_INIT=16'b1100011101100101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI767P1_0_9_LC_4_13_5  (
            .in0(N__16399),
            .in1(N__16168),
            .in2(N__16704),
            .in3(N__20474),
            .lcout(),
            .ltout(\this_vga_signals.N_24_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_4_13_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_4_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__16162),
            .in2(N__16102),
            .in3(N__16098),
            .lcout(),
            .ltout(\this_vga_signals.g0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_4_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_4_13_7 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_LC_4_13_7  (
            .in0(N__16075),
            .in1(N__16060),
            .in2(N__16030),
            .in3(N__16027),
            .lcout(\this_vga_signals.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_8_LC_4_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_8_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3SF72_8_LC_4_14_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3SF72_8_LC_4_14_0  (
            .in0(N__18849),
            .in1(N__15994),
            .in2(N__16450),
            .in3(N__19091),
            .lcout(\this_vga_signals.g0_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_4_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_4_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI13H13_9_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__20025),
            .in2(_gnd_net_),
            .in3(N__19880),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI13H13Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_4_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_4_15_3 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_4_15_3  (
            .in0(N__16213),
            .in1(N__15982),
            .in2(N__19099),
            .in3(N__18937),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_16_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_16_6  (
            .in0(N__17146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16997),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_8_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_8_0 .LUT_INIT=16'b1001101001011001;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_0_LC_5_8_0  (
            .in0(N__16889),
            .in1(N__18127),
            .in2(N__18526),
            .in3(N__17704),
            .lcout(),
            .ltout(\this_vga_signals.if_N_8_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_8_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_8_1 .LUT_INIT=16'b0011000011110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_1_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__18622),
            .in2(N__16201),
            .in3(N__18375),
            .lcout(),
            .ltout(\this_vga_signals.if_N_9_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_5_8_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_5_8_2 .LUT_INIT=16'b0100011100011101;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_0_LC_5_8_2  (
            .in0(N__18623),
            .in1(N__18507),
            .in2(N__16198),
            .in3(N__18441),
            .lcout(\this_vga_signals.mult1_un82_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_8_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_8_5 .LUT_INIT=16'b1100100110010011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_0_LC_5_8_5  (
            .in0(N__17705),
            .in1(N__16890),
            .in2(N__18527),
            .in3(N__18128),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_5_9_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_5_9_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIVC6I_0_LC_5_9_0  (
            .in0(N__18317),
            .in1(N__18364),
            .in2(N__18329),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_d7lt4 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_5_9_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_5_9_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_5_9_1  (
            .in0(N__20072),
            .in1(N__18640),
            .in2(_gnd_net_),
            .in3(N__16195),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_3_LC_5_9_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_5_9_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_5_9_2  (
            .in0(N__20065),
            .in1(N__18523),
            .in2(_gnd_net_),
            .in3(N__16192),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_4_LC_5_9_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_5_9_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_5_9_3  (
            .in0(N__20073),
            .in1(N__18129),
            .in2(_gnd_net_),
            .in3(N__16189),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_5_LC_5_9_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_5_9_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_5_9_4  (
            .in0(N__20066),
            .in1(N__18197),
            .in2(_gnd_net_),
            .in3(N__16186),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_6_LC_5_9_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_5_9_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_5_9_5  (
            .in0(N__20074),
            .in1(N__19001),
            .in2(_gnd_net_),
            .in3(N__16429),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_7_LC_5_9_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_5_9_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_5_9_6  (
            .in0(N__20067),
            .in1(N__19069),
            .in2(_gnd_net_),
            .in3(N__16426),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_8_LC_5_9_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_5_9_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_5_9_7  (
            .in0(N__20075),
            .in1(N__18819),
            .in2(_gnd_net_),
            .in3(N__16423),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__40354),
            .ce(),
            .sr(N__16516));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_5_10_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_5_10_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__18924),
            .in2(_gnd_net_),
            .in3(N__16420),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40367),
            .ce(N__16477),
            .sr(N__16514));
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m5_i_a4_0_0_LC_5_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_m5_i_a4_0_0_LC_5_11_1  (
            .in0(N__18534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18400),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclto3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_5_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_5_11_2 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIADGD1_5_LC_5_11_2  (
            .in0(N__18644),
            .in1(N__18209),
            .in2(N__16417),
            .in3(N__18140),
            .lcout(\this_vga_signals.un4_hsynclto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_d_0_sqmuxa_1_0_o2_LC_5_11_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_d_0_sqmuxa_1_0_o2_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_d_0_sqmuxa_1_0_o2_LC_5_11_5 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \this_ppu.M_vaddress_d_0_sqmuxa_1_0_o2_LC_5_11_5  (
            .in0(N__16414),
            .in1(N__16687),
            .in2(_gnd_net_),
            .in3(N__16400),
            .lcout(\this_ppu.N_759_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_5_12_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16324),
            .lcout(this_vga_signals_M_vcounter_q_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40387),
            .ce(N__16300),
            .sr(N__16257));
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_8_LC_5_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_8_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNISKQ82_8_LC_5_13_1 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNISKQ82_8_LC_5_13_1  (
            .in0(N__19092),
            .in1(N__16222),
            .in2(N__18853),
            .in3(N__19014),
            .lcout(\this_vga_signals.un4_hsynclt9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_5_13_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_2_LC_5_13_7 .LUT_INIT=16'b1001110001100011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_2_LC_5_13_7  (
            .in0(N__16818),
            .in1(N__16681),
            .in2(N__17597),
            .in3(N__17343),
            .lcout(\this_vga_signals.g0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_1_LC_5_14_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_1_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_1_LC_5_14_0 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_1_LC_5_14_0  (
            .in0(N__16609),
            .in1(N__17344),
            .in2(_gnd_net_),
            .in3(N__16602),
            .lcout(\this_vga_signals.g0_0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_5_14_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_5_14_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_5_14_2  (
            .in0(N__16495),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20029),
            .lcout(\this_vga_signals.N_935_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_5_14_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_5_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16462),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40409),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_5_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_5_14_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIGR3I_9_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__18928),
            .in2(_gnd_net_),
            .in3(N__20478),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_0_9_LC_5_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_0_9_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_0_9_LC_5_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIQJSA2_0_9_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19718),
            .lcout(M_vcounter_q_esr_RNIQJSA2_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_5_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_5_6 .LUT_INIT=16'b0101000001011010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_6_5_6  (
            .in0(N__17841),
            .in1(_gnd_net_),
            .in2(N__17901),
            .in3(N__17952),
            .lcout(\this_vga_ramdac.N_24_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_6_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_6_7 .LUT_INIT=16'b0101011101010011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_6_6_7  (
            .in0(N__17995),
            .in1(N__17960),
            .in2(N__17852),
            .in3(N__17897),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_7_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_7_4 .LUT_INIT=16'b0100101100010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_6_7_4  (
            .in0(N__17892),
            .in1(N__17853),
            .in2(N__17962),
            .in3(N__17997),
            .lcout(\this_vga_ramdac.m16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_7_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_7_5 .LUT_INIT=16'b0101100100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_6_7_5  (
            .in0(N__17998),
            .in1(N__17842),
            .in2(N__17961),
            .in3(N__17891),
            .lcout(\this_vga_ramdac.m19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_6_7_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_6_7_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_0_0_LC_6_7_6  (
            .in0(N__18571),
            .in1(N__17671),
            .in2(N__17041),
            .in3(N__18444),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_7_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_7_7 .LUT_INIT=16'b0001010100111101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_6_7_7  (
            .in0(N__17996),
            .in1(N__17956),
            .in2(N__17857),
            .in3(N__17893),
            .lcout(\this_vga_ramdac.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIFBB7K_1_LC_6_8_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIFBB7K_1_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIFBB7K_1_LC_6_8_1 .LUT_INIT=16'b1100001100111010;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIFBB7K_1_LC_6_8_1  (
            .in0(N__18624),
            .in1(N__18383),
            .in2(N__18528),
            .in3(N__18427),
            .lcout(),
            .ltout(\this_vga_signals.d_N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_am_LC_6_8_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_am_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_am_LC_6_8_2 .LUT_INIT=16'b1001000011110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_am_LC_6_8_2  (
            .in0(N__18384),
            .in1(N__18625),
            .in2(N__17032),
            .in3(N__17733),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_2_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_8_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_8_3 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_8_3  (
            .in0(N__17029),
            .in1(N__17650),
            .in2(N__17019),
            .in3(N__23973),
            .lcout(\this_vga_ramdac.N_2687_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_9_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_6_9_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_6_9_0  (
            .in0(N__17646),
            .in1(N__18049),
            .in2(N__16959),
            .in3(N__23956),
            .lcout(\this_vga_ramdac.N_28_i_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_9_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_9_2 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_6_9_2  (
            .in0(N__17645),
            .in1(N__16924),
            .in2(N__16908),
            .in3(N__23955),
            .lcout(\this_vga_ramdac.N_2690_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_9_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_9_3 .LUT_INIT=16'b1000100110011101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_LC_6_9_3  (
            .in0(N__16891),
            .in1(N__18116),
            .in2(N__18525),
            .in3(N__17706),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_9_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_LC_6_9_4  (
            .in0(N__17707),
            .in1(N__18064),
            .in2(N__16873),
            .in3(N__18268),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_6_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_6_9_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_2_LC_6_9_5  (
            .in0(N__18607),
            .in1(N__17152),
            .in2(N__18524),
            .in3(N__18115),
            .lcout(\this_vga_signals.M_hcounter_d7lt7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_6_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_6_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc1_LC_6_9_7  (
            .in0(N__18500),
            .in1(N__18117),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_10_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_10_0 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_6_10_0  (
            .in0(N__17644),
            .in1(N__17803),
            .in2(N__17139),
            .in3(N__23960),
            .lcout(\this_vga_ramdac.N_2691_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40355),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_6_10_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_LC_6_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__19159),
            .in2(_gnd_net_),
            .in3(N__18282),
            .lcout(\this_vga_signals.pixel_clk_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40355),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_10_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_10_2 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_6_10_2  (
            .in0(N__17643),
            .in1(N__17122),
            .in2(N__17106),
            .in3(N__23959),
            .lcout(\this_vga_ramdac.N_2689_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40355),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_6_10_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_6_10_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI6MKH3_4_LC_6_10_3  (
            .in0(N__17089),
            .in1(N__17080),
            .in2(_gnd_net_),
            .in3(N__17599),
            .lcout(\this_vga_signals.N_819_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_6_10_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_6_10_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIF4AR_5_LC_6_10_4  (
            .in0(N__18196),
            .in1(N__19053),
            .in2(_gnd_net_),
            .in3(N__18997),
            .lcout(\this_vga_signals.M_lcounter_q_3_i_o2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI4VLK7_LC_6_10_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI4VLK7_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNI4VLK7_LC_6_10_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNI4VLK7_LC_6_10_5  (
            .in0(N__19179),
            .in1(N__19158),
            .in2(_gnd_net_),
            .in3(N__18281),
            .lcout(M_pcounter_q_ret_1_RNI4VLK7),
            .ltout(M_pcounter_q_ret_1_RNI4VLK7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_10_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_10_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_6_10_6  (
            .in0(N__17052),
            .in1(N__17071),
            .in2(N__17062),
            .in3(N__23957),
            .lcout(\this_vga_ramdac.N_2686_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40355),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_10_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_10_7 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_6_10_7  (
            .in0(N__23958),
            .in1(N__17659),
            .in2(N__17616),
            .in3(N__17642),
            .lcout(\this_vga_ramdac.N_2688_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40355),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_6_11_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_1_LC_6_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_1_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__17584),
            .in2(_gnd_net_),
            .in3(N__17391),
            .lcout(\this_vga_signals.g0_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_6_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_0_LC_6_11_2 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_0_LC_6_11_2  (
            .in0(N__19134),
            .in1(N__20057),
            .in2(N__19183),
            .in3(N__19849),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40368),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_6_15_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_6_15_2 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_6_15_2  (
            .in0(N__19098),
            .in1(N__18936),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(M_hcounter_q_esr_RNIU8TO_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI63POP1_9_LC_7_4_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI63POP1_9_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI63POP1_9_LC_7_4_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI63POP1_9_LC_7_4_0  (
            .in0(N__17773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18057),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UV2O8_9_LC_7_4_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UV2O8_9_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4UV2O8_9_LC_7_4_1 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI4UV2O8_9_LC_7_4_1  (
            .in0(N__17752),
            .in1(N__17179),
            .in2(N__18058),
            .in3(N__17782),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4GRFM_9_LC_7_4_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4GRFM_9_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4GRFM_9_LC_7_4_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI4GRFM_9_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(N__18051),
            .in2(_gnd_net_),
            .in3(N__18448),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI50QR8_9_LC_7_4_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI50QR8_9_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI50QR8_9_LC_7_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI50QR8_9_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__18056),
            .in2(_gnd_net_),
            .in3(N__17719),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4T6U44_9_LC_7_4_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4T6U44_9_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI4T6U44_9_LC_7_4_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI4T6U44_9_LC_7_4_7  (
            .in0(N__18052),
            .in1(N__17178),
            .in2(_gnd_net_),
            .in3(N__17772),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7U1Q5_9_LC_7_5_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7U1Q5_9_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI7U1Q5_9_LC_7_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI7U1Q5_9_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__18220),
            .in2(_gnd_net_),
            .in3(N__18050),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_7_6_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_7_6_4 .LUT_INIT=16'b0100001001110101;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_7_6_4  (
            .in0(N__17994),
            .in1(N__17943),
            .in2(N__17902),
            .in3(N__17846),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_7_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_7_1 .LUT_INIT=16'b1101001010110100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_7_7_1  (
            .in0(N__18570),
            .in1(N__17670),
            .in2(N__17743),
            .in3(N__18443),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_7_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m5_i_LC_7_7_3 .LUT_INIT=16'b0010011001100100;
    LogicCell40 \this_vga_signals.un4_haddress_if_m5_i_LC_7_7_3  (
            .in0(N__18646),
            .in1(N__18397),
            .in2(N__18547),
            .in3(N__18442),
            .lcout(),
            .ltout(\this_vga_signals.N_2_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.haddress_1_0_LC_7_7_4 .C_ON=1'b0;
    defparam \this_vga_signals.haddress_1_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.haddress_1_0_LC_7_7_4 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \this_vga_signals.haddress_1_0_LC_7_7_4  (
            .in0(N__17677),
            .in1(N__17765),
            .in2(N__17791),
            .in3(N__17788),
            .lcout(\this_vga_signals.haddress_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_7_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_7_5 .LUT_INIT=16'b0010000101111011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_m2_LC_7_7_5  (
            .in0(N__17766),
            .in1(N__18398),
            .in2(N__18654),
            .in3(N__18292),
            .lcout(\this_vga_signals.mult1_un89_sum_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_bm_LC_7_7_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_bm_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_bm_LC_7_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_2_bm_LC_7_7_7  (
            .in0(N__17739),
            .in1(N__18141),
            .in2(_gnd_net_),
            .in3(N__17715),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_2_bm ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_8_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_8_4 .LUT_INIT=16'b0010001010111011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_c2_LC_7_8_4  (
            .in0(N__18542),
            .in1(N__18645),
            .in2(_gnd_net_),
            .in3(N__18428),
            .lcout(\this_vga_signals.mult1_un75_sum_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_7_8_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_x4_LC_7_8_6 .LUT_INIT=16'b1001001100110110;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_x4_LC_7_8_6  (
            .in0(N__18650),
            .in1(N__18563),
            .in2(N__18546),
            .in3(N__18429),
            .lcout(),
            .ltout(\this_vga_signals.if_N_8_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_8_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_8_7 .LUT_INIT=16'b0011000011110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__18399),
            .in2(N__18334),
            .in3(N__18330),
            .lcout(\this_vga_signals.if_N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_7_9_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_7_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18283),
            .lcout(\this_vga_signals.M_pcounter_q_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40334),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_7_9_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_7_9_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNIB85C3_LC_7_9_4  (
            .in0(N__19135),
            .in1(N__19146),
            .in2(_gnd_net_),
            .in3(N__19839),
            .lcout(),
            .ltout(\this_vga_signals.M_pcounter_q_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_1_LC_7_9_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_1_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_1_LC_7_9_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNIR5V44_1_LC_7_9_5  (
            .in0(N__20006),
            .in1(_gnd_net_),
            .in2(N__18286),
            .in3(N__19108),
            .lcout(\this_vga_signals.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_7_9_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_7_9_6 .LUT_INIT=16'b1100111010001100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_c3_LC_7_9_6  (
            .in0(N__18267),
            .in1(N__18238),
            .in2(N__18211),
            .in3(N__19008),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_7_9_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_7_9_7 .LUT_INIT=16'b0110010110100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_axbxc3_1_0_LC_7_9_7  (
            .in0(N__19009),
            .in1(N__18208),
            .in2(N__18145),
            .in3(N__18133),
            .lcout(\this_vga_signals.mult1_un68_sum_axbxc3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOSP33_9_LC_7_10_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOSP33_9_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIOSP33_9_LC_7_10_2 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIOSP33_9_LC_7_10_2  (
            .in0(N__18920),
            .in1(N__18840),
            .in2(N__19710),
            .in3(N__19097),
            .lcout(N_28_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_7_10_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_7_10_6 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIC8KO2_9_LC_7_10_6  (
            .in0(N__18019),
            .in1(N__18919),
            .in2(N__19192),
            .in3(N__18839),
            .lcout(\this_vga_signals.N_83_1 ),
            .ltout(\this_vga_signals.N_83_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIGO4F3_LC_7_10_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIGO4F3_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_1_RNIGO4F3_LC_7_10_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_1_RNIGO4F3_LC_7_10_7  (
            .in0(N__20030),
            .in1(N__19178),
            .in2(N__19162),
            .in3(N__19132),
            .lcout(\this_vga_signals.N_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_7_11_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_1_LC_7_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_1_LC_7_11_2  (
            .in0(N__19150),
            .in1(N__19133),
            .in2(_gnd_net_),
            .in3(N__19848),
            .lcout(\this_vga_signals.M_pcounter_q_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40356),
            .ce(N__20063),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_7_12_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_7_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIBP6I_7_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__19096),
            .in2(_gnd_net_),
            .in3(N__19015),
            .lcout(),
            .ltout(\this_vga_signals.N_809_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT8TC3_9_LC_7_12_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT8TC3_9_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIT8TC3_9_LC_7_12_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIT8TC3_9_LC_7_12_6  (
            .in0(N__19711),
            .in1(N__18932),
            .in2(N__18856),
            .in3(N__18847),
            .lcout(N_34_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5I298_9_LC_7_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5I298_9_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI5I298_9_LC_7_16_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI5I298_9_LC_7_16_2  (
            .in0(N__29229),
            .in1(N__37753),
            .in2(_gnd_net_),
            .in3(N__19719),
            .lcout(port_nmib_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_9_21_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_9_21_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_9_21_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_0_LC_9_21_0 (
            .in0(N__22858),
            .in1(N__18729),
            .in2(N__22160),
            .in3(N__22136),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_1_LC_9_21_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_9_21_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_9_21_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_1_LC_9_21_1 (
            .in0(N__22864),
            .in1(N__18702),
            .in2(_gnd_net_),
            .in3(N__18688),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_2_LC_9_21_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_9_21_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_9_21_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_2_LC_9_21_2 (
            .in0(N__22859),
            .in1(N__18672),
            .in2(_gnd_net_),
            .in3(N__18658),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_3_LC_9_21_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_9_21_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_9_21_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_3_LC_9_21_3 (
            .in0(N__22865),
            .in1(N__19398),
            .in2(_gnd_net_),
            .in3(N__19384),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_4_LC_9_21_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_9_21_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_9_21_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_4_LC_9_21_4 (
            .in0(N__22860),
            .in1(N__19368),
            .in2(_gnd_net_),
            .in3(N__19354),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_5_LC_9_21_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_9_21_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_9_21_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_5_LC_9_21_5 (
            .in0(N__22862),
            .in1(N__19341),
            .in2(_gnd_net_),
            .in3(N__19327),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_6_LC_9_21_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_9_21_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_9_21_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_6_LC_9_21_6 (
            .in0(N__22861),
            .in1(N__19314),
            .in2(_gnd_net_),
            .in3(N__19300),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_7_LC_9_21_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_9_21_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_9_21_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_7_LC_9_21_7 (
            .in0(N__22863),
            .in1(N__19284),
            .in2(_gnd_net_),
            .in3(N__19270),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__40436),
            .ce(),
            .sr(N__28898));
    defparam M_this_map_address_q_8_LC_9_22_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_9_22_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_9_22_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_8_LC_9_22_0 (
            .in0(N__22866),
            .in1(N__19254),
            .in2(_gnd_net_),
            .in3(N__19240),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__40444),
            .ce(),
            .sr(N__28896));
    defparam M_this_map_address_q_9_LC_9_22_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_9_22_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_9_22_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_map_address_q_9_LC_9_22_1 (
            .in0(N__19224),
            .in1(N__22867),
            .in2(_gnd_net_),
            .in3(N__19237),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40444),
            .ce(),
            .sr(N__28896));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_10_8_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_10_8_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI67JU6_9_LC_10_8_2  (
            .in0(N__20024),
            .in1(N__19870),
            .in2(N__19449),
            .in3(N__20512),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNI67JU6Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_10_14_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_10_14_7 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_10_14_7  (
            .in0(N__19445),
            .in1(N__19881),
            .in2(N__20608),
            .in3(N__20513),
            .lcout(\this_vga_signals.N_826_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_10_16_5 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_10_16_5 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_10_16_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_10_16_5  (
            .in0(N__19666),
            .in1(N__19794),
            .in2(_gnd_net_),
            .in3(N__39882),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40371),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_406_LC_10_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.G_406_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_406_LC_10_16_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.G_406_LC_10_16_7  (
            .in0(N__19665),
            .in1(N__19793),
            .in2(_gnd_net_),
            .in3(N__39881),
            .lcout(\this_vga_signals.GZ0Z_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_0_LC_10_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_0_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_0_LC_10_20_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_0_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__35608),
            .in2(_gnd_net_),
            .in3(N__22162),
            .lcout(M_this_map_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_3_LC_10_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_3_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_3_LC_10_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_3_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__39517),
            .in2(_gnd_net_),
            .in3(N__22135),
            .lcout(M_this_map_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_4_LC_10_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_4_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_4_LC_10_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_4_LC_10_23_1  (
            .in0(N__41039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22173),
            .lcout(M_this_map_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI8K9F5_0_1_LC_11_10_3.C_ON=1'b0;
    defparam M_this_state_q_RNI8K9F5_0_1_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI8K9F5_0_1_LC_11_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 M_this_state_q_RNI8K9F5_0_1_LC_11_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29225),
            .lcout(dma_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_14_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_14_5 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_14_5  (
            .in0(N__19450),
            .in1(N__19892),
            .in2(N__20552),
            .in3(N__20514),
            .lcout(),
            .ltout(\this_vga_signals.N_827_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_11_14_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_11_14_6 .LUT_INIT=16'b0111010011001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_11_14_6  (
            .in0(N__19893),
            .in1(N__20607),
            .in2(N__19417),
            .in3(N__19987),
            .lcout(this_vga_signals_M_lcounter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40336),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_11_15_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_11_15_3 .LUT_INIT=16'b0011100011111000;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_11_15_3  (
            .in0(N__19414),
            .in1(N__19955),
            .in2(N__20554),
            .in3(N__19891),
            .lcout(this_vga_signals_M_lcounter_q_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40345),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_11_16_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_11_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19795),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40358),
            .ce(),
            .sr(N__39784));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_1_LC_11_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_1_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_1_LC_11_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_1_LC_11_20_3  (
            .in0(_gnd_net_),
            .in1(N__35504),
            .in2(_gnd_net_),
            .in3(N__22161),
            .lcout(M_this_map_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_2_LC_11_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_2_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_2_LC_11_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_2_LC_11_21_4  (
            .in0(N__22163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38764),
            .lcout(M_this_map_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_7_LC_11_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_7_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_7_LC_11_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_7_LC_11_23_4  (
            .in0(N__22165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36478),
            .lcout(M_this_map_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_5_LC_11_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_5_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_5_LC_11_23_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_5_LC_11_23_6  (
            .in0(N__22164),
            .in1(N__40608),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_map_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIAJH46_5_LC_12_9_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIAJH46_5_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIAJH46_5_LC_12_9_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIAJH46_5_LC_12_9_3  (
            .in0(N__21529),
            .in1(N__24174),
            .in2(N__31642),
            .in3(N__21646),
            .lcout(M_this_ppu_vram_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIITCPC_LC_12_11_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIITCPC_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIITCPC_LC_12_11_0 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIITCPC_LC_12_11_0  (
            .in0(N__19720),
            .in1(N__23954),
            .in2(N__29224),
            .in3(N__29982),
            .lcout(\this_ppu.M_last_q_RNIITCPC ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_0_LC_12_12_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_0_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_0_LC_12_12_4 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \this_ppu.M_vaddress_q_0_LC_12_12_4  (
            .in0(N__24085),
            .in1(N__29148),
            .in2(N__31843),
            .in3(N__24031),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40312),
            .ce(),
            .sr(N__29756));
    defparam \this_ppu.line_clk.M_last_q_LC_12_14_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_12_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_12_14_3  (
            .in0(N__20606),
            .in1(N__20581),
            .in2(N__20553),
            .in3(N__20518),
            .lcout(\this_ppu.M_last_q ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40327),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_srsts_0_i_o2_1_0_LC_12_15_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_srsts_0_i_o2_1_0_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_srsts_0_i_o2_1_0_LC_12_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_srsts_0_i_o2_1_0_LC_12_15_5  (
            .in0(N__20602),
            .in1(N__20580),
            .in2(N__20551),
            .in3(N__20511),
            .lcout(\this_ppu.N_5_4 ),
            .ltout(\this_ppu.N_5_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_12_15_6 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_12_15_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_12_15_6  (
            .in0(N__24066),
            .in1(_gnd_net_),
            .in2(N__20404),
            .in3(N__29141),
            .lcout(\this_ppu.N_228_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_0_LC_12_21_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_0_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_0_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_0_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20401),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40400),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_12_21_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_12_21_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_12_21_4  (
            .in0(N__20383),
            .in1(N__34923),
            .in2(_gnd_net_),
            .in3(N__20377),
            .lcout(M_this_ppu_spr_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_1_LC_12_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_1_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_1_LC_12_22_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_1_LC_12_22_1  (
            .in0(N__31862),
            .in1(N__31790),
            .in2(_gnd_net_),
            .in3(N__29968),
            .lcout(\this_ppu.M_vaddress_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40410),
            .ce(),
            .sr(N__29769));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_13_7_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_13_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_13_7_4  (
            .in0(N__38914),
            .in1(N__20137),
            .in2(_gnd_net_),
            .in3(N__20122),
            .lcout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIQER3C_9_LC_13_8_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIQER3C_9_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIQER3C_9_LC_13_8_3 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \this_ppu.M_state_q_RNIQER3C_9_LC_13_8_3  (
            .in0(N__29640),
            .in1(N__24769),
            .in2(_gnd_net_),
            .in3(N__29560),
            .lcout(M_state_q_RNIQER3C_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI1IH46_4_LC_13_9_0 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI1IH46_4_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI1IH46_4_LC_13_9_0 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNI1IH46_4_LC_13_9_0  (
            .in0(N__24172),
            .in1(N__21527),
            .in2(N__31687),
            .in3(N__21853),
            .lcout(M_this_ppu_vram_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIBKH46_6_LC_13_9_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIBKH46_6_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIBKH46_6_LC_13_9_2 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIBKH46_6_LC_13_9_2  (
            .in0(N__24173),
            .in1(N__21528),
            .in2(N__31594),
            .in3(N__21991),
            .lcout(M_this_ppu_vram_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNI0B6K1_3_LC_13_9_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNI0B6K1_3_LC_13_9_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNI0B6K1_3_LC_13_9_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNI0B6K1_3_LC_13_9_7  (
            .in0(N__28277),
            .in1(N__31734),
            .in2(_gnd_net_),
            .in3(N__24171),
            .lcout(\this_ppu.N_806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIF0FG4_3_LC_13_10_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIF0FG4_3_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIF0FG4_3_LC_13_10_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIF0FG4_3_LC_13_10_3  (
            .in0(N__28278),
            .in1(N__24178),
            .in2(N__31738),
            .in3(N__21556),
            .lcout(M_this_ppu_vram_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_11_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_11_6  (
            .in0(N__38901),
            .in1(N__21499),
            .in2(_gnd_net_),
            .in3(N__21484),
            .lcout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_18_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_18_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_13_18_3  (
            .in0(N__21715),
            .in1(N__21469),
            .in2(_gnd_net_),
            .in3(N__34975),
            .lcout(M_this_ppu_spr_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_20_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_13_20_0  (
            .in0(N__27985),
            .in1(N__21256),
            .in2(_gnd_net_),
            .in3(N__34956),
            .lcout(M_this_ppu_spr_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_20_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_20_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_20_4  (
            .in0(N__20614),
            .in1(N__21049),
            .in2(_gnd_net_),
            .in3(N__34957),
            .lcout(M_this_ppu_spr_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_20_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_20_6  (
            .in0(N__29692),
            .in1(N__20857),
            .in2(_gnd_net_),
            .in3(N__34958),
            .lcout(M_this_ppu_spr_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_3_LC_13_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_3_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20629),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40391),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_2_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21730),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40391),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_6_LC_13_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_6_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_ram_write_data_0_a2_6_LC_13_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_map_ram_write_data_0_a2_6_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(N__36278),
            .in2(_gnd_net_),
            .in3(N__22166),
            .lcout(M_this_map_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_14_8_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_14_8_1 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_14_8_1  (
            .in0(N__22262),
            .in1(N__21598),
            .in2(N__22327),
            .in3(N__21697),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_14_9_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_14_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_LC_14_9_4  (
            .in0(N__21691),
            .in1(N__21670),
            .in2(_gnd_net_),
            .in3(N__38935),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_14_9_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_14_9_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_14_9_5  (
            .in0(N__22264),
            .in1(N__38980),
            .in2(N__21655),
            .in3(N__21652),
            .lcout(M_this_spr_ram_read_data_2),
            .ltout(M_this_spr_ram_read_data_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vram_en_0_i_o2_LC_14_9_6 .C_ON=1'b0;
    defparam \this_ppu.vram_en_0_i_o2_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vram_en_0_i_o2_LC_14_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.vram_en_0_i_o2_LC_14_9_6  (
            .in0(N__21990),
            .in1(N__21849),
            .in2(N__21637),
            .in3(N__21555),
            .lcout(\this_ppu.N_772_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_14_9_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_14_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_14_9_7  (
            .in0(N__38934),
            .in1(N__21634),
            .in2(_gnd_net_),
            .in3(N__21616),
            .lcout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_14_10_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_14_10_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_14_10_3  (
            .in0(N__21592),
            .in1(N__21574),
            .in2(_gnd_net_),
            .in3(N__38943),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_14_10_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_14_10_4 .LUT_INIT=16'b1011100100110001;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_14_10_4  (
            .in0(N__22263),
            .in1(N__21748),
            .in2(N__21559),
            .in3(N__38812),
            .lcout(M_this_spr_ram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_14_10_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_14_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_14_10_6  (
            .in0(N__38944),
            .in1(N__21826),
            .in2(_gnd_net_),
            .in3(N__21808),
            .lcout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_14_11_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_14_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_14_11_0  (
            .in0(N__38933),
            .in1(N__21793),
            .in2(_gnd_net_),
            .in3(N__21775),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_14_11_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_14_11_1 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_14_11_1  (
            .in0(N__22323),
            .in1(N__22247),
            .in2(N__21757),
            .in3(N__21754),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_3_LC_14_12_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_3_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_3_LC_14_12_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_3_LC_14_12_0  (
            .in0(N__28275),
            .in1(N__28380),
            .in2(_gnd_net_),
            .in3(N__21909),
            .lcout(M_this_ppu_vram_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40305),
            .ce(),
            .sr(N__22414));
    defparam \this_delay_clk.M_pipe_q_2_LC_14_14_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21742),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40313),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_1_LC_14_18_1.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_14_18_1.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_14_18_1.LUT_INIT=16'b0000011000001100;
    LogicCell40 M_this_oam_address_q_1_LC_14_18_1 (
            .in0(N__24602),
            .in1(N__24698),
            .in2(N__25018),
            .in3(N__24655),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40346),
            .ce(),
            .sr(N__28895));
    defparam \this_ppu.M_state_q_8_LC_14_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_8_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_8_LC_14_19_2 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \this_ppu.M_state_q_8_LC_14_19_2  (
            .in0(N__24133),
            .in1(N__24757),
            .in2(N__28552),
            .in3(N__29580),
            .lcout(\this_ppu.M_state_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40359),
            .ce(),
            .sr(N__39777));
    defparam M_this_oam_address_q_RNI24IA1_1_LC_14_20_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_14_20_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_14_20_4.LUT_INIT=16'b1111111100100000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_LC_14_20_4 (
            .in0(N__24701),
            .in1(N__24657),
            .in2(N__24603),
            .in3(N__39883),
            .lcout(N_1286_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_14_21_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_14_21_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_14_21_7.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_0_1_LC_14_21_7 (
            .in0(N__24702),
            .in1(N__24658),
            .in2(N__24604),
            .in3(N__39891),
            .lcout(N_1294_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_6_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_6_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_6_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_15_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_15_9_6 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_15_9_6  (
            .in0(N__21859),
            .in1(N__36127),
            .in2(N__22261),
            .in3(N__22030),
            .lcout(M_this_spr_ram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNI1O64C_1_LC_15_10_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNI1O64C_1_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNI1O64C_1_LC_15_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_ppu.M_haddress_q_RNI1O64C_1_LC_15_10_0  (
            .in0(N__27938),
            .in1(N__29330),
            .in2(N__28356),
            .in3(N__21928),
            .lcout(\this_ppu.un1_M_haddress_q_c3 ),
            .ltout(\this_ppu.un1_M_haddress_q_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_RNIHAI4C_5_LC_15_10_1 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIHAI4C_5_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIHAI4C_5_LC_15_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_haddress_q_RNIHAI4C_5_LC_15_10_1  (
            .in0(N__28194),
            .in1(N__28117),
            .in2(N__21838),
            .in3(N__28285),
            .lcout(\this_ppu.un1_M_haddress_q_c6 ),
            .ltout(\this_ppu.un1_M_haddress_q_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_6_LC_15_10_2 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_6_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_6_LC_15_10_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_ppu.M_haddress_q_6_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21835),
            .in3(N__28067),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40291),
            .ce(),
            .sr(N__22409));
    defparam \this_ppu.M_state_q_RNIQER3C_0_9_LC_15_10_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIQER3C_0_9_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIQER3C_0_9_LC_15_10_3 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \this_ppu.M_state_q_RNIQER3C_0_9_LC_15_10_3  (
            .in0(N__29632),
            .in1(N__24765),
            .in2(_gnd_net_),
            .in3(N__29556),
            .lcout(\this_ppu.N_754_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_5_LC_15_10_7 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_5_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_5_LC_15_10_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_haddress_q_5_LC_15_10_7  (
            .in0(N__28195),
            .in1(N__28118),
            .in2(N__28295),
            .in3(N__21832),
            .lcout(M_this_ppu_vram_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40291),
            .ce(),
            .sr(N__22409));
    defparam \this_ppu.M_haddress_q_RNIJU24C_1_LC_15_11_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_RNIJU24C_1_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_haddress_q_RNIJU24C_1_LC_15_11_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_haddress_q_RNIJU24C_1_LC_15_11_5  (
            .in0(N__27942),
            .in1(N__29319),
            .in2(_gnd_net_),
            .in3(N__21929),
            .lcout(\this_ppu.un1_M_haddress_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_15_11_7 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_15_11_7 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_15_11_7  (
            .in0(N__29139),
            .in1(N__24038),
            .in2(N__24099),
            .in3(N__39894),
            .lcout(\this_ppu.M_last_q_RNIGL6V4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_4_LC_15_12_0 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_4_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_4_LC_15_12_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \this_ppu.M_haddress_q_4_LC_15_12_0  (
            .in0(N__28276),
            .in1(N__28347),
            .in2(N__28196),
            .in3(N__21910),
            .lcout(M_this_ppu_vram_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40300),
            .ce(),
            .sr(N__22405));
    defparam M_this_oam_address_q_0_LC_15_15_1.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_15_15_1.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_15_15_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_0_LC_15_15_1 (
            .in0(N__25006),
            .in1(N__24582),
            .in2(_gnd_net_),
            .in3(N__24643),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40314),
            .ce(),
            .sr(N__28897));
    defparam \this_ppu.M_state_q_9_LC_15_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_9_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_9_LC_15_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.M_state_q_9_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21898),
            .lcout(\this_ppu.M_state_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40347),
            .ce(),
            .sr(N__39774));
    defparam M_this_data_tmp_q_esr_13_LC_15_21_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_15_21_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_15_21_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_15_21_1 (
            .in0(N__40600),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40372),
            .ce(N__29039),
            .sr(N__39781));
    defparam \this_ppu.M_state_q_0_LC_15_22_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_15_22_4 .SEQ_MODE=4'b1001;
    defparam \this_ppu.M_state_q_0_LC_15_22_4 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \this_ppu.M_state_q_0_LC_15_22_4  (
            .in0(N__29115),
            .in1(N__23115),
            .in2(N__24103),
            .in3(N__24043),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40380),
            .ce(),
            .sr(N__39785));
    defparam \this_ppu.M_count_q_7_LC_15_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_7_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_7_LC_15_22_7 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_ppu.M_count_q_7_LC_15_22_7  (
            .in0(N__23114),
            .in1(N__22504),
            .in2(_gnd_net_),
            .in3(N__30010),
            .lcout(\this_ppu.M_count_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40380),
            .ce(),
            .sr(N__39785));
    defparam \this_ppu.M_state_q_RNINUC91_4_LC_15_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNINUC91_4_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNINUC91_4_LC_15_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNINUC91_4_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__29448),
            .in2(_gnd_net_),
            .in3(N__29670),
            .lcout(\this_ppu.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_10_LC_15_24_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_15_24_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_15_24_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_15_24_0 (
            .in0(N__38769),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40401),
            .ce(N__29046),
            .sr(N__39793));
    defparam M_this_data_tmp_q_esr_12_LC_15_25_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_15_25_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_15_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_15_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41054),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40411),
            .ce(N__29057),
            .sr(N__39794));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_16_8_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_16_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_16_8_4  (
            .in0(N__38932),
            .in1(N__21892),
            .in2(_gnd_net_),
            .in3(N__21877),
            .lcout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_16_9_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_16_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_16_9_2  (
            .in0(N__38931),
            .in1(N__22066),
            .in2(_gnd_net_),
            .in3(N__22051),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_16_9_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_16_9_3 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_16_9_3  (
            .in0(N__22318),
            .in1(N__22233),
            .in2(N__22033),
            .in3(N__21943),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_16_9_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_16_9_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_spr_ram.mem_mem_4_0_wclke_3_LC_16_9_4  (
            .in0(N__37549),
            .in1(N__37374),
            .in2(N__37477),
            .in3(N__37300),
            .lcout(\this_spr_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_16_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_16_9_6 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_12_LC_16_9_6  (
            .in0(N__22234),
            .in1(N__22000),
            .in2(N__22567),
            .in3(N__22319),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_16_9_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_16_9_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_11_LC_16_9_7  (
            .in0(N__22254),
            .in1(N__22525),
            .in2(N__21994),
            .in3(N__33550),
            .lcout(M_this_spr_ram_read_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_16_10_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_16_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_16_10_7  (
            .in0(N__38930),
            .in1(N__21973),
            .in2(_gnd_net_),
            .in3(N__21958),
            .lcout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_haddress_q_7_LC_16_11_3 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_7_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_7_LC_16_11_3 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \this_ppu.M_haddress_q_7_LC_16_11_3  (
            .in0(N__28032),
            .in1(N__28066),
            .in2(_gnd_net_),
            .in3(N__21937),
            .lcout(\this_ppu.M_haddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40290),
            .ce(),
            .sr(N__22413));
    defparam \this_ppu.M_haddress_q_2_LC_16_11_4 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_2_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_2_LC_16_11_4 .LUT_INIT=16'b1001110011001100;
    LogicCell40 \this_ppu.M_haddress_q_2_LC_16_11_4  (
            .in0(N__21931),
            .in1(N__28375),
            .in2(N__29338),
            .in3(N__27944),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40290),
            .ce(),
            .sr(N__22413));
    defparam \this_ppu.M_haddress_q_1_LC_16_11_5 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_1_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_1_LC_16_11_5 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \this_ppu.M_haddress_q_1_LC_16_11_5  (
            .in0(N__27943),
            .in1(N__29323),
            .in2(_gnd_net_),
            .in3(N__21930),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40290),
            .ce(),
            .sr(N__22413));
    defparam \this_ppu.M_haddress_q_0_LC_16_11_6 .C_ON=1'b0;
    defparam \this_ppu.M_haddress_q_0_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_haddress_q_0_LC_16_11_6 .LUT_INIT=16'b0101101000011110;
    LogicCell40 \this_ppu.M_haddress_q_0_LC_16_11_6  (
            .in0(N__29641),
            .in1(N__24764),
            .in2(N__29337),
            .in3(N__29579),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40290),
            .ce(),
            .sr(N__22413));
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_16_12_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_16_12_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_wclke_3_LC_16_12_2  (
            .in0(N__37358),
            .in1(N__37304),
            .in2(N__37462),
            .in3(N__37529),
            .lcout(\this_spr_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_12_LC_16_12_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_12_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_12_LC_16_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_12_LC_16_12_3  (
            .in0(N__28969),
            .in1(N__22348),
            .in2(_gnd_net_),
            .in3(N__34976),
            .lcout(\this_spr_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40295),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_0 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_16_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22291),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40304),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_11_LC_16_15_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_11_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_11_LC_16_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_radreg_11_LC_16_15_3  (
            .in0(N__22282),
            .in1(N__22975),
            .in2(_gnd_net_),
            .in3(N__34962),
            .lcout(\this_spr_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40308),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_a2_LC_16_17_4 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_a2_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_a2_LC_16_17_4 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \this_ppu.un1_M_this_state_q_1_i_0_0_a2_LC_16_17_4  (
            .in0(N__24454),
            .in1(N__36739),
            .in2(N__24487),
            .in3(N__24530),
            .lcout(M_this_state_d_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_16_18_7.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_16_18_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_3_LC_16_18_7 (
            .in0(N__23026),
            .in1(N__24903),
            .in2(_gnd_net_),
            .in3(N__23046),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40326),
            .ce(N__24815),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_16_19_0.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_16_19_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_16_19_0.LUT_INIT=16'b0100111001000100;
    LogicCell40 M_this_data_count_q_10_LC_16_19_0 (
            .in0(N__24909),
            .in1(N__23809),
            .in2(N__39922),
            .in3(N__22827),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40335),
            .ce(N__24823),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_11_LC_16_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_11_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_6_11_LC_16_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_6_11_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__23047),
            .in2(_gnd_net_),
            .in3(N__23069),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_6Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_16_19_3.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_16_19_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_16_19_3.LUT_INIT=16'b0000000010100101;
    LogicCell40 M_this_data_count_q_11_LC_16_19_3 (
            .in0(N__23796),
            .in1(_gnd_net_),
            .in2(N__23782),
            .in3(N__24904),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40335),
            .ce(N__24823),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_11_LC_16_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_11_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_7_11_LC_16_19_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_7_11_LC_16_19_4  (
            .in0(N__23219),
            .in1(N__23795),
            .in2(N__24937),
            .in3(N__23820),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_i_a2_7Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_11_LC_16_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_11_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_11_LC_16_19_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_11_LC_16_19_5  (
            .in0(N__23101),
            .in1(N__23128),
            .in2(N__22429),
            .in3(N__22426),
            .lcout(\this_ppu.N_934 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_16_19_6.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_16_19_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_16_19_6.LUT_INIT=16'b0000101000000101;
    LogicCell40 M_this_data_count_q_12_LC_16_19_6 (
            .in0(N__23220),
            .in1(_gnd_net_),
            .in2(N__24910),
            .in3(N__23206),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40335),
            .ce(N__24823),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_16_19_7.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_16_19_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_16_19_7.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_2_LC_16_19_7 (
            .in0(N__23056),
            .in1(N__24908),
            .in2(_gnd_net_),
            .in3(N__23070),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40335),
            .ce(N__24823),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_6_LC_16_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_6_LC_16_20_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_6_LC_16_20_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_ppu.M_state_q_6_LC_16_20_0  (
            .in0(_gnd_net_),
            .in1(N__28545),
            .in2(_gnd_net_),
            .in3(N__24126),
            .lcout(\this_ppu.M_state_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40344),
            .ce(),
            .sr(N__39775));
    defparam M_this_data_tmp_q_esr_20_LC_16_21_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_16_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_16_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_16_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41055),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40357),
            .ce(N__32422),
            .sr(N__39778));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_22_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_c_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(N__25039),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_22_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_0_s1_THRU_LUT4_0_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__23874),
            .in2(N__23768),
            .in3(N__22420),
            .lcout(\this_ppu.un1_M_count_q_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_0_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_22_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_1_s1_THRU_LUT4_0_LC_16_22_2  (
            .in0(_gnd_net_),
            .in1(N__23759),
            .in2(N__22489),
            .in3(N__22417),
            .lcout(\this_ppu.un1_M_count_q_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_1_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_22_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_2_s1_THRU_LUT4_0_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(N__22617),
            .in2(N__23769),
            .in3(N__22519),
            .lcout(\this_ppu.un1_M_count_q_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_2_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_22_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_3_s1_THRU_LUT4_0_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(N__23763),
            .in2(N__22452),
            .in3(N__22516),
            .lcout(\this_ppu.un1_M_count_q_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_3_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_22_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_4_s1_THRU_LUT4_0_LC_16_22_5  (
            .in0(_gnd_net_),
            .in1(N__23991),
            .in2(N__23770),
            .in3(N__22513),
            .lcout(\this_ppu.un1_M_count_q_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_4_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_22_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_count_q_1_cry_5_s1_THRU_LUT4_0_LC_16_22_6  (
            .in0(_gnd_net_),
            .in1(N__23767),
            .in2(N__22645),
            .in3(N__22510),
            .lcout(\this_ppu.un1_M_count_q_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_count_q_1_cry_5_s1 ),
            .carryout(\this_ppu.un1_M_count_q_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNO_0_7_LC_16_22_7 .LUT_INIT=16'b1100110000110110;
    LogicCell40 \this_ppu.M_count_q_RNO_0_7_LC_16_22_7  (
            .in0(N__29449),
            .in1(N__23857),
            .in2(N__30022),
            .in3(N__22507),
            .lcout(\this_ppu.M_count_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_2_LC_16_23_0 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_2_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_2_LC_16_23_0 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_2_LC_16_23_0  (
            .in0(N__22488),
            .in1(N__25093),
            .in2(N__22498),
            .in3(N__25063),
            .lcout(\this_ppu.M_count_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40379),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIDE0G_2_LC_16_23_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_count_q_RNIDE0G_2_LC_16_23_2  (
            .in0(N__23990),
            .in1(N__22445),
            .in2(N__22644),
            .in3(N__22484),
            .lcout(),
            .ltout(\this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIKM001_1_LC_16_23_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.M_count_q_RNIKM001_1_LC_16_23_3  (
            .in0(N__22613),
            .in1(N__23873),
            .in2(N__22468),
            .in3(N__23842),
            .lcout(\this_ppu.M_hoffset_d_0_sqmuxa_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_4_LC_16_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_4_LC_16_23_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_4_LC_16_23_4 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_4_LC_16_23_4  (
            .in0(N__22453),
            .in1(N__25094),
            .in2(N__22465),
            .in3(N__25065),
            .lcout(\this_ppu.M_count_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40379),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_6_LC_16_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_6_LC_16_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_6_LC_16_23_5 .LUT_INIT=16'b1010100000000010;
    LogicCell40 \this_ppu.M_count_q_6_LC_16_23_5  (
            .in0(N__25066),
            .in1(N__25096),
            .in2(N__22654),
            .in3(N__22640),
            .lcout(\this_ppu.M_count_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40379),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_3_LC_16_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_3_LC_16_23_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_3_LC_16_23_7 .LUT_INIT=16'b1010000010000010;
    LogicCell40 \this_ppu.M_count_q_3_LC_16_23_7  (
            .in0(N__25064),
            .in1(N__25095),
            .in2(N__22618),
            .in3(N__22624),
            .lcout(\this_ppu.M_count_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40379),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_16_LC_16_24_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_16_24_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_16_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_16_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35588),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40390),
            .ce(N__32423),
            .sr(N__39790));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_31_5.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_31_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_31_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_16_31_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39889),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_17_9_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_17_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_17_9_0  (
            .in0(N__38936),
            .in1(N__22591),
            .in2(_gnd_net_),
            .in3(N__22579),
            .lcout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_17_9_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_17_9_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_17_9_1  (
            .in0(N__24234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22558),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40287),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_17_9_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_17_9_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_17_9_4  (
            .in0(N__24187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24233),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40287),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_17_9_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_17_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_17_9_7  (
            .in0(N__22552),
            .in1(N__22540),
            .in2(_gnd_net_),
            .in3(N__38937),
            .lcout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_17_10_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_17_10_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__24255),
            .in2(_gnd_net_),
            .in3(N__22792),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40292),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_6_LC_17_10_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_17_10_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__24258),
            .in2(_gnd_net_),
            .in3(N__22810),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40292),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_17_10_6 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_17_10_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_17_10_6  (
            .in0(N__24257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22798),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40292),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_17_10_7 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_17_10_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__24256),
            .in2(_gnd_net_),
            .in3(N__22804),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40292),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_17_11_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_17_11_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_17_11_2  (
            .in0(N__24260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22786),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40296),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_17_11_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_17_11_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__22780),
            .in2(_gnd_net_),
            .in3(N__24259),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40296),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_17_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_17_12_0  (
            .in0(N__24261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40301),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_17_14_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_17_14_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__22774),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40309),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_17_14_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_17_14_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_spr_ram.mem_mem_2_0_wclke_3_LC_17_14_3  (
            .in0(N__37341),
            .in1(N__37273),
            .in2(N__37441),
            .in3(N__37500),
            .lcout(\this_spr_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_17_14_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_17_14_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_2_LC_17_14_4  (
            .in0(N__38791),
            .in1(N__37193),
            .in2(N__36294),
            .in3(N__36657),
            .lcout(M_this_spr_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_5_LC_17_15_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_5_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_5_LC_17_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_5_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22993),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40315),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_17_15_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_17_15_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \this_start_data_delay.M_last_q_LC_17_15_6  (
            .in0(N__24531),
            .in1(N__24449),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(this_start_data_delay_M_last_q),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40315),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_17_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_17_16_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_1_LC_17_16_2  (
            .in0(N__35511),
            .in1(N__37183),
            .in2(N__40609),
            .in3(N__36678),
            .lcout(M_this_spr_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_10_LC_17_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_10_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_10_LC_17_16_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_10_LC_17_16_4  (
            .in0(N__24477),
            .in1(N__24511),
            .in2(_gnd_net_),
            .in3(N__24450),
            .lcout(\this_ppu.N_321_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_map_address_q_0_i_o2_0_a2_4_LC_17_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_map_address_q_0_i_o2_0_a2_4_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_map_address_q_0_i_o2_0_a2_4_LC_17_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_map_address_q_0_i_o2_0_a2_4_LC_17_16_6  (
            .in0(N__30577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40803),
            .lcout(N_609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_17_17_2.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_17_17_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_17_17_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_4_LC_17_17_2 (
            .in0(N__23017),
            .in1(N__24900),
            .in2(_gnd_net_),
            .in3(N__23147),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40328),
            .ce(N__24819),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_17_17_3.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_17_17_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_17_17_3.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_5_LC_17_17_3 (
            .in0(N__24901),
            .in1(N__23008),
            .in2(_gnd_net_),
            .in3(N__23193),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40328),
            .ce(N__24819),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_17_17_4.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_17_17_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_17_17_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_9_LC_17_17_4 (
            .in0(N__23833),
            .in1(N__24902),
            .in2(_gnd_net_),
            .in3(N__23168),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40328),
            .ce(N__24819),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_17_17_6.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_17_17_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_17_17_6.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_0_LC_17_17_6 (
            .in0(N__23091),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24899),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40328),
            .ce(N__24819),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_11_LC_17_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_11_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_9_11_LC_17_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_9_11_LC_17_17_7  (
            .in0(N__24387),
            .in1(N__24410),
            .in2(N__24357),
            .in3(N__23090),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_9Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_c_0_LC_17_18_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_17_18_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_17_18_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_17_18_0 (
            .in0(_gnd_net_),
            .in1(N__23092),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_17_18_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_17_18_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_17_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_17_18_1 (
            .in0(_gnd_net_),
            .in1(N__24411),
            .in2(N__23694),
            .in3(N__23077),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_17_18_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_17_18_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_17_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_17_18_2 (
            .in0(_gnd_net_),
            .in1(N__23640),
            .in2(N__23074),
            .in3(N__23050),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_17_18_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_17_18_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_17_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_17_18_3 (
            .in0(_gnd_net_),
            .in1(N__23045),
            .in2(N__23695),
            .in3(N__23020),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_17_18_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_17_18_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_17_18_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_17_18_4 (
            .in0(_gnd_net_),
            .in1(N__23644),
            .in2(N__23152),
            .in3(N__23011),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_17_18_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_17_18_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_17_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_17_18_5 (
            .in0(_gnd_net_),
            .in1(N__23192),
            .in2(N__23696),
            .in3(N__23002),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_17_18_6.C_ON=1'b1;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_17_18_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_17_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_5_THRU_LUT4_0_LC_17_18_6 (
            .in0(_gnd_net_),
            .in1(N__23648),
            .in2(N__24388),
            .in3(N__22999),
            .lcout(M_this_data_count_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_17_18_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_17_18_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_17_18_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_17_18_7 (
            .in0(_gnd_net_),
            .in1(N__23697),
            .in2(N__24358),
            .in3(N__22996),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_17_19_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_17_19_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_17_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_17_19_0 (
            .in0(_gnd_net_),
            .in1(N__24835),
            .in2(N__23755),
            .in3(N__23836),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_17_19_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_17_19_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_17_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_8_THRU_LUT4_0_LC_17_19_1 (
            .in0(_gnd_net_),
            .in1(N__23172),
            .in2(N__23749),
            .in3(N__23824),
            .lcout(M_this_data_count_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_10_LC_17_19_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_10_LC_17_19_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_10_LC_17_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_10_LC_17_19_2 (
            .in0(_gnd_net_),
            .in1(N__23821),
            .in2(N__23754),
            .in3(N__23803),
            .lcout(M_this_data_count_q_s_10),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_17_19_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_17_19_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_17_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_10_THRU_LUT4_0_LC_17_19_3 (
            .in0(_gnd_net_),
            .in1(N__23735),
            .in2(N__23800),
            .in3(N__23773),
            .lcout(M_this_data_count_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_17_19_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_17_19_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_17_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_11_THRU_LUT4_0_LC_17_19_4 (
            .in0(_gnd_net_),
            .in1(N__23708),
            .in2(N__23224),
            .in3(N__23200),
            .lcout(M_this_data_count_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_13_LC_17_19_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_13_LC_17_19_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_13_LC_17_19_5.LUT_INIT=16'b1010101001010101;
    LogicCell40 M_this_data_count_q_RNO_0_13_LC_17_19_5 (
            .in0(N__24933),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23197),
            .lcout(M_this_data_count_q_s_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_11_LC_17_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_11_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_a2_8_11_LC_17_19_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_a2_8_11_LC_17_19_6  (
            .in0(N__24834),
            .in1(N__23194),
            .in2(N__23173),
            .in3(N__23148),
            .lcout(\this_ppu.M_this_state_q_srsts_i_a2_8Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_17_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_17_20_6 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \this_ppu.M_state_q_5_LC_17_20_6  (
            .in0(N__28511),
            .in1(N__23122),
            .in2(N__29455),
            .in3(N__29734),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40360),
            .ce(),
            .sr(N__39772));
    defparam \this_ppu.M_state_q_RNIEOOI_9_LC_17_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIEOOI_9_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIEOOI_9_LC_17_21_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_state_q_RNIEOOI_9_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__29625),
            .in2(_gnd_net_),
            .in3(N__24729),
            .lcout(\this_ppu.N_760_0 ),
            .ltout(\this_ppu.N_760_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIKDTE1_5_LC_17_21_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIKDTE1_5_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIKDTE1_5_LC_17_21_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_state_q_RNIKDTE1_5_LC_17_21_3  (
            .in0(N__24124),
            .in1(N__29520),
            .in2(N__24181),
            .in3(N__41436),
            .lcout(\this_ppu.N_762_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII6H51_5_LC_17_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII6H51_5_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII6H51_5_LC_17_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNII6H51_5_LC_17_21_5  (
            .in0(N__24730),
            .in1(N__24125),
            .in2(N__29447),
            .in3(N__28507),
            .lcout(\this_ppu.M_state_q_inv_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI7O615_LC_17_22_0 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI7O615_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI7O615_LC_17_22_0 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI7O615_LC_17_22_0  (
            .in0(N__24098),
            .in1(N__29443),
            .in2(N__29140),
            .in3(N__24039),
            .lcout(\this_ppu.N_268_i_0_0 ),
            .ltout(\this_ppu.N_268_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_5_LC_17_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_5_LC_17_22_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_5_LC_17_22_1 .LUT_INIT=16'b1010100100000000;
    LogicCell40 \this_ppu.M_count_q_5_LC_17_22_1  (
            .in0(N__23992),
            .in1(N__24001),
            .in2(N__23995),
            .in3(N__25062),
            .lcout(\this_ppu.M_count_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40381),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI7KJ86_0_4_LC_17_22_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI7KJ86_0_4_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI7KJ86_0_4_LC_17_22_3 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_ppu.M_state_q_RNI7KJ86_0_4_LC_17_22_3  (
            .in0(N__29674),
            .in1(N__23953),
            .in2(N__29451),
            .in3(N__29983),
            .lcout(\this_ppu.N_1323_0 ),
            .ltout(\this_ppu.N_1323_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_1_LC_17_22_4 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_1_LC_17_22_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_1_LC_17_22_4 .LUT_INIT=16'b1100000010010000;
    LogicCell40 \this_ppu.M_count_q_1_LC_17_22_4  (
            .in0(N__23887),
            .in1(N__23875),
            .in2(N__23878),
            .in3(N__25092),
            .lcout(\this_ppu.M_count_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40381),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_count_q_RNIL508_7_LC_17_22_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_count_q_RNIL508_7_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__23856),
            .in2(_gnd_net_),
            .in3(N__25034),
            .lcout(\this_ppu.M_hoffset_d_0_sqmuxa_0_a3_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_6_LC_17_23_5.C_ON=1'b0;
    defparam M_this_oam_address_q_6_LC_17_23_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_6_LC_17_23_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_6_LC_17_23_5 (
            .in0(N__24317),
            .in1(N__25011),
            .in2(_gnd_net_),
            .in3(N__25107),
            .lcout(M_this_oam_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40392),
            .ce(),
            .sr(N__28891));
    defparam M_this_oam_address_q_7_LC_17_24_2.C_ON=1'b0;
    defparam M_this_oam_address_q_7_LC_17_24_2.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_7_LC_17_24_2.LUT_INIT=16'b0001001000110000;
    LogicCell40 M_this_oam_address_q_7_LC_17_24_2 (
            .in0(N__24318),
            .in1(N__25013),
            .in2(N__24285),
            .in3(N__25108),
            .lcout(M_this_oam_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40402),
            .ce(),
            .sr(N__28890));
    defparam M_this_oam_address_q_2_LC_17_24_3.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_17_24_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_17_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_oam_address_q_2_LC_17_24_3 (
            .in0(N__25012),
            .in1(N__25295),
            .in2(_gnd_net_),
            .in3(N__25227),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40402),
            .ce(),
            .sr(N__28890));
    defparam M_this_data_tmp_q_esr_9_LC_17_25_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_17_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_17_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_17_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35491),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40412),
            .ce(N__29053),
            .sr(N__39791));
    defparam M_this_data_tmp_q_esr_18_LC_17_27_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_17_27_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_17_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_17_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38780),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40426),
            .ce(N__32427),
            .sr(N__39795));
    defparam \this_reset_cond.M_stage_q_7_LC_18_10_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_18_10_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_18_10_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_18_10_0  (
            .in0(N__24262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24193),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40297),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_13_LC_18_13_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_13_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_13_LC_18_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_13_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__32183),
            .in2(_gnd_net_),
            .in3(N__30634),
            .lcout(\this_ppu.N_324_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_18_14_5.C_ON=1'b0;
    defparam M_this_state_q_9_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_18_14_5.LUT_INIT=16'b0000000010001000;
    LogicCell40 M_this_state_q_9_LC_18_14_5 (
            .in0(N__40805),
            .in1(N__28950),
            .in2(_gnd_net_),
            .in3(N__39913),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_7_LC_18_14_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_7_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_7_LC_18_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_7_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__30547),
            .in2(_gnd_net_),
            .in3(N__40804),
            .lcout(N_332_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_en_1_sqmuxa_0_a2_i_o2_LC_18_15_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_en_1_sqmuxa_0_a2_i_o2_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_en_1_sqmuxa_0_a2_i_o2_LC_18_15_0 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_en_1_sqmuxa_0_a2_i_o2_LC_18_15_0  (
            .in0(N__36799),
            .in1(N__24475),
            .in2(N__24541),
            .in3(N__24442),
            .lcout(N_314_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.N_660_i_LC_18_15_1 .C_ON=1'b0;
    defparam \this_ppu.N_660_i_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.N_660_i_LC_18_15_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \this_ppu.N_660_i_LC_18_15_1  (
            .in0(N__24476),
            .in1(N__30625),
            .in2(_gnd_net_),
            .in3(N__39897),
            .lcout(N_660_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_address_q_0_i_o3_0_a2_0_LC_18_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_address_q_0_i_o3_0_a2_0_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_address_q_0_i_o3_0_a2_0_LC_18_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_address_q_0_i_o3_0_a2_0_LC_18_15_2  (
            .in0(N__32310),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40819),
            .lcout(N_611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_18_15_5.C_ON=1'b0;
    defparam M_this_state_q_8_LC_18_15_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_18_15_5.LUT_INIT=16'b1100110010000000;
    LogicCell40 M_this_state_q_8_LC_18_15_5 (
            .in0(N__30329),
            .in1(N__32136),
            .in2(N__32275),
            .in3(N__28948),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40321),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_18_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_18_15_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_12_LC_18_15_6  (
            .in0(N__24540),
            .in1(N__24474),
            .in2(_gnd_net_),
            .in3(N__24441),
            .lcout(N_309_0),
            .ltout(N_309_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_LC_18_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_LC_18_15_7 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_LC_18_15_7  (
            .in0(_gnd_net_),
            .in1(N__28947),
            .in2(N__24421),
            .in3(N__36656),
            .lcout(N_260_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_qlde_0_i_i_LC_18_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_qlde_0_i_i_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_qlde_0_i_i_LC_18_16_0 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \this_ppu.M_this_data_count_qlde_0_i_i_LC_18_16_0  (
            .in0(N__40794),
            .in1(N__30664),
            .in2(N__40664),
            .in3(N__39890),
            .lcout(N_257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_1_0_LC_18_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_1_0_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_a2_1_0_LC_18_16_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_a2_1_0_LC_18_16_5  (
            .in0(N__28949),
            .in1(N__36677),
            .in2(_gnd_net_),
            .in3(N__40793),
            .lcout(\this_ppu.N_545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_18_17_0.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_18_17_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_18_17_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_1_LC_18_17_0 (
            .in0(N__24418),
            .in1(N__24873),
            .in2(_gnd_net_),
            .in3(N__24412),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40337),
            .ce(N__24811),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_18_17_2.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_18_17_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_18_17_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_6_LC_18_17_2 (
            .in0(N__24394),
            .in1(N__24874),
            .in2(_gnd_net_),
            .in3(N__24386),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40337),
            .ce(N__24811),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_18_17_3.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_18_17_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_18_17_3.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_7_LC_18_17_3 (
            .in0(N__24875),
            .in1(N__24364),
            .in2(_gnd_net_),
            .in3(N__24356),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40337),
            .ce(N__24811),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_18_17_5.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_18_17_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_18_17_5.LUT_INIT=16'b0101000011011000;
    LogicCell40 M_this_data_count_q_13_LC_18_17_5 (
            .in0(N__24876),
            .in1(N__30450),
            .in2(N__24949),
            .in3(N__39914),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40337),
            .ce(N__24811),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a2_0_a2_LC_18_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a2_0_a2_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a2_0_a2_LC_18_18_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_sqmuxa_0_a2_0_a2_LC_18_18_3  (
            .in0(N__24645),
            .in1(N__24571),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(M_this_oam_ram_write_data_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIMU531_1_LC_18_18_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIMU531_1_LC_18_18_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIMU531_1_LC_18_18_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIMU531_1_LC_18_18_7 (
            .in0(N__24644),
            .in1(N__24699),
            .in2(N__36811),
            .in3(N__40836),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_18_19_5.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_18_19_5.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_18_19_5.LUT_INIT=16'b0010001011100010;
    LogicCell40 M_this_data_count_q_8_LC_18_19_5 (
            .in0(N__24916),
            .in1(N__24898),
            .in2(N__25014),
            .in3(N__39915),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40361),
            .ce(N__24804),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_7_LC_18_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_7_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_7_LC_18_20_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_7_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__28515),
            .in2(_gnd_net_),
            .in3(N__29730),
            .lcout(\this_ppu.M_state_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40373),
            .ce(),
            .sr(N__39767));
    defparam \this_ppu.M_oamcurr_q_3_LC_18_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_3_LC_18_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_3_LC_18_21_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oamcurr_q_3_LC_18_21_4  (
            .in0(N__30168),
            .in1(N__28437),
            .in2(_gnd_net_),
            .in3(N__28806),
            .lcout(M_this_ppu_oam_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40382),
            .ce(),
            .sr(N__28893));
    defparam \this_ppu.M_oamcurr_q_RNIRKBD7_4_LC_18_22_4 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNIRKBD7_4_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNIRKBD7_4_LC_18_22_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNIRKBD7_4_LC_18_22_4  (
            .in0(N__30164),
            .in1(N__25366),
            .in2(_gnd_net_),
            .in3(N__28804),
            .lcout(\this_ppu.un1_M_oamcurr_q_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIRE716_4_LC_18_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIRE716_4_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIRE716_4_LC_18_22_5 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \this_ppu.M_state_q_RNIRE716_4_LC_18_22_5  (
            .in0(N__29450),
            .in1(N__29683),
            .in2(_gnd_net_),
            .in3(N__30000),
            .lcout(\this_ppu.M_oamcurr_qc_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_18_22_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_18_22_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_18_22_6.LUT_INIT=16'b1111111100010000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_1_LC_18_22_6 (
            .in0(N__24706),
            .in1(N__24656),
            .in2(N__24595),
            .in3(N__39896),
            .lcout(N_1302_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_count_q_0_LC_18_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_count_q_0_LC_18_22_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_count_q_0_LC_18_22_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \this_ppu.M_count_q_0_LC_18_22_7  (
            .in0(N__25038),
            .in1(N__25091),
            .in2(_gnd_net_),
            .in3(N__25061),
            .lcout(\this_ppu.M_count_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40393),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_3_LC_18_23_0.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_18_23_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_18_23_0.LUT_INIT=16'b0001010001010000;
    LogicCell40 M_this_oam_address_q_3_LC_18_23_0 (
            .in0(N__24993),
            .in1(N__25296),
            .in2(N__25254),
            .in3(N__25228),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_1_LC_18_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_1_LC_18_23_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_1_LC_18_23_1 .LUT_INIT=16'b1100000001001000;
    LogicCell40 \this_ppu.M_oamcurr_q_1_LC_18_23_1  (
            .in0(N__28736),
            .in1(N__28435),
            .in2(N__28674),
            .in3(N__28621),
            .lcout(M_this_ppu_oam_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam M_this_oam_address_q_4_LC_18_23_2.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_18_23_2.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_18_23_2.LUT_INIT=16'b0000010100001010;
    LogicCell40 M_this_oam_address_q_4_LC_18_23_2 (
            .in0(N__25203),
            .in1(_gnd_net_),
            .in2(N__25010),
            .in3(N__25130),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam M_this_oam_address_q_5_LC_18_23_3.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_18_23_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_18_23_3.LUT_INIT=16'b0001001000110000;
    LogicCell40 M_this_oam_address_q_5_LC_18_23_3 (
            .in0(N__25131),
            .in1(N__24994),
            .in2(N__25179),
            .in3(N__25204),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_4_LC_18_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_4_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_4_LC_18_23_4 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_oamcurr_q_4_LC_18_23_4  (
            .in0(N__28436),
            .in1(N__25367),
            .in2(N__30183),
            .in3(N__28807),
            .lcout(M_this_ppu_oam_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_0_LC_18_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_0_LC_18_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_0_LC_18_23_5 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \this_ppu.M_oamcurr_q_0_LC_18_23_5  (
            .in0(N__28735),
            .in1(N__28432),
            .in2(_gnd_net_),
            .in3(N__28620),
            .lcout(M_this_ppu_oam_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_5_LC_18_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_5_LC_18_23_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_5_LC_18_23_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \this_ppu.M_oamcurr_q_5_LC_18_23_6  (
            .in0(N__28434),
            .in1(N__28463),
            .in2(_gnd_net_),
            .in3(N__28407),
            .lcout(M_this_ppu_oam_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_2_LC_18_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_2_LC_18_23_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_2_LC_18_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_oamcurr_q_2_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(N__28433),
            .in2(_gnd_net_),
            .in3(N__28840),
            .lcout(M_this_ppu_oam_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40403),
            .ce(),
            .sr(N__28892));
    defparam \this_ppu.M_oamcurr_q_RNI3AD1_4_LC_18_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNI3AD1_4_LC_18_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNI3AD1_4_LC_18_24_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_oamcurr_q_RNI3AD1_4_LC_18_24_2  (
            .in0(N__30066),
            .in1(N__28657),
            .in2(N__25377),
            .in3(N__28727),
            .lcout(\this_ppu.M_state_q_srsts_i_i_o2_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_1_LC_18_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_1_LC_18_24_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamidx_q_1_LC_18_24_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oamidx_q_1_LC_18_24_3  (
            .in0(N__30286),
            .in1(N__39912),
            .in2(N__30259),
            .in3(N__30020),
            .lcout(\this_ppu.M_oamidx_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40413),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_13_LC_18_24_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_13_LC_18_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_13_LC_18_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_13_LC_18_24_5  (
            .in0(N__25339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39269),
            .lcout(M_this_oam_ram_write_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNILNG41_3_LC_18_24_6.C_ON=1'b0;
    defparam M_this_oam_address_q_RNILNG41_3_LC_18_24_6.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNILNG41_3_LC_18_24_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNILNG41_3_LC_18_24_6 (
            .in0(N__25294),
            .in1(N__25247),
            .in2(_gnd_net_),
            .in3(N__25220),
            .lcout(un1_M_this_oam_address_q_c4),
            .ltout(un1_M_this_oam_address_q_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIOKR51_5_LC_18_24_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_18_24_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_18_24_7.LUT_INIT=16'b1010000000000000;
    LogicCell40 M_this_oam_address_q_RNIOKR51_5_LC_18_24_7 (
            .in0(N__25178),
            .in1(_gnd_net_),
            .in2(N__25153),
            .in3(N__25129),
            .lcout(un1_M_this_oam_address_q_c6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_8_LC_18_25_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_18_25_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_18_25_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_18_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35602),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40420),
            .ce(N__29065),
            .sr(N__39786));
    defparam M_this_data_tmp_q_esr_15_LC_18_25_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_18_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_18_25_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_18_25_4 (
            .in0(N__36472),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40420),
            .ce(N__29065),
            .sr(N__39786));
    defparam M_this_data_tmp_q_esr_11_LC_18_25_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_18_25_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_18_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_18_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39498),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40420),
            .ce(N__29065),
            .sr(N__39786));
    defparam M_this_data_tmp_q_esr_21_LC_18_26_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_18_26_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_18_26_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_18_26_0 (
            .in0(N__40598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40427),
            .ce(N__32438),
            .sr(N__39792));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_18_LC_18_27_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_18_LC_18_27_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_18_LC_18_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_18_LC_18_27_2  (
            .in0(_gnd_net_),
            .in1(N__27001),
            .in2(_gnd_net_),
            .in3(N__39270),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_21_LC_18_27_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_21_LC_18_27_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_21_LC_18_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_21_LC_18_27_4  (
            .in0(_gnd_net_),
            .in1(N__26980),
            .in2(_gnd_net_),
            .in3(N__39271),
            .lcout(M_this_oam_ram_write_data_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_spr_address_q_0_LC_19_13_0.C_ON=1'b1;
    defparam M_this_spr_address_q_0_LC_19_13_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_0_LC_19_13_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_0_LC_19_13_0 (
            .in0(N__30442),
            .in1(N__26772),
            .in2(N__28921),
            .in3(N__28920),
            .lcout(M_this_spr_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_19_13_0_),
            .carryout(un1_M_this_spr_address_q_cry_0),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_1_LC_19_13_1.C_ON=1'b1;
    defparam M_this_spr_address_q_1_LC_19_13_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_1_LC_19_13_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_1_LC_19_13_1 (
            .in0(N__30446),
            .in1(N__26576),
            .in2(_gnd_net_),
            .in3(N__26527),
            .lcout(M_this_spr_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_0),
            .carryout(un1_M_this_spr_address_q_cry_1),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_2_LC_19_13_2.C_ON=1'b1;
    defparam M_this_spr_address_q_2_LC_19_13_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_2_LC_19_13_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_2_LC_19_13_2 (
            .in0(N__30443),
            .in1(N__26340),
            .in2(_gnd_net_),
            .in3(N__26320),
            .lcout(M_this_spr_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_1),
            .carryout(un1_M_this_spr_address_q_cry_2),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_3_LC_19_13_3.C_ON=1'b1;
    defparam M_this_spr_address_q_3_LC_19_13_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_3_LC_19_13_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_3_LC_19_13_3 (
            .in0(N__30447),
            .in1(N__26090),
            .in2(_gnd_net_),
            .in3(N__26065),
            .lcout(M_this_spr_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_2),
            .carryout(un1_M_this_spr_address_q_cry_3),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_4_LC_19_13_4.C_ON=1'b1;
    defparam M_this_spr_address_q_4_LC_19_13_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_4_LC_19_13_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_4_LC_19_13_4 (
            .in0(N__30444),
            .in1(N__25889),
            .in2(_gnd_net_),
            .in3(N__25876),
            .lcout(M_this_spr_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_3),
            .carryout(un1_M_this_spr_address_q_cry_4),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_5_LC_19_13_5.C_ON=1'b1;
    defparam M_this_spr_address_q_5_LC_19_13_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_5_LC_19_13_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_5_LC_19_13_5 (
            .in0(N__30448),
            .in1(N__25687),
            .in2(_gnd_net_),
            .in3(N__25648),
            .lcout(M_this_spr_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_4),
            .carryout(un1_M_this_spr_address_q_cry_5),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_6_LC_19_13_6.C_ON=1'b1;
    defparam M_this_spr_address_q_6_LC_19_13_6.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_6_LC_19_13_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_6_LC_19_13_6 (
            .in0(N__30445),
            .in1(N__25407),
            .in2(_gnd_net_),
            .in3(N__25387),
            .lcout(M_this_spr_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_5),
            .carryout(un1_M_this_spr_address_q_cry_6),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_7_LC_19_13_7.C_ON=1'b1;
    defparam M_this_spr_address_q_7_LC_19_13_7.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_7_LC_19_13_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_7_LC_19_13_7 (
            .in0(N__30449),
            .in1(N__27695),
            .in2(_gnd_net_),
            .in3(N__27670),
            .lcout(M_this_spr_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_6),
            .carryout(un1_M_this_spr_address_q_cry_7),
            .clk(N__40317),
            .ce(),
            .sr(N__28900));
    defparam M_this_spr_address_q_8_LC_19_14_0.C_ON=1'b1;
    defparam M_this_spr_address_q_8_LC_19_14_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_8_LC_19_14_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_8_LC_19_14_0 (
            .in0(N__30414),
            .in1(N__27484),
            .in2(_gnd_net_),
            .in3(N__27457),
            .lcout(M_this_spr_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_19_14_0_),
            .carryout(un1_M_this_spr_address_q_cry_8),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_spr_address_q_9_LC_19_14_1.C_ON=1'b1;
    defparam M_this_spr_address_q_9_LC_19_14_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_9_LC_19_14_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_9_LC_19_14_1 (
            .in0(N__30417),
            .in1(N__27267),
            .in2(_gnd_net_),
            .in3(N__27250),
            .lcout(M_this_spr_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_8),
            .carryout(un1_M_this_spr_address_q_cry_9),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_spr_address_q_10_LC_19_14_2.C_ON=1'b1;
    defparam M_this_spr_address_q_10_LC_19_14_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_10_LC_19_14_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_10_LC_19_14_2 (
            .in0(N__30412),
            .in1(N__27052),
            .in2(_gnd_net_),
            .in3(N__27013),
            .lcout(M_this_spr_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_9),
            .carryout(un1_M_this_spr_address_q_cry_10),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_spr_address_q_11_LC_19_14_3.C_ON=1'b1;
    defparam M_this_spr_address_q_11_LC_19_14_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_11_LC_19_14_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_11_LC_19_14_3 (
            .in0(N__30416),
            .in1(N__37260),
            .in2(_gnd_net_),
            .in3(N__27010),
            .lcout(M_this_spr_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_10),
            .carryout(un1_M_this_spr_address_q_cry_11),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_spr_address_q_12_LC_19_14_4.C_ON=1'b1;
    defparam M_this_spr_address_q_12_LC_19_14_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_12_LC_19_14_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_12_LC_19_14_4 (
            .in0(N__30413),
            .in1(N__37340),
            .in2(_gnd_net_),
            .in3(N__27007),
            .lcout(M_this_spr_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_11),
            .carryout(un1_M_this_spr_address_q_cry_12),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_spr_address_q_13_LC_19_14_5.C_ON=1'b0;
    defparam M_this_spr_address_q_13_LC_19_14_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_13_LC_19_14_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_spr_address_q_13_LC_19_14_5 (
            .in0(N__37421),
            .in1(N__30415),
            .in2(_gnd_net_),
            .in3(N__27004),
            .lcout(M_this_spr_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40322),
            .ce(),
            .sr(N__28899));
    defparam M_this_state_q_RNILR691_2_LC_19_15_2.C_ON=1'b0;
    defparam M_this_state_q_RNILR691_2_LC_19_15_2.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNILR691_2_LC_19_15_2.LUT_INIT=16'b1111111110001000;
    LogicCell40 M_this_state_q_RNILR691_2_LC_19_15_2 (
            .in0(N__32602),
            .in1(N__40827),
            .in2(_gnd_net_),
            .in3(N__39903),
            .lcout(N_1310_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_12_LC_19_15_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_12_LC_19_15_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_12_LC_19_15_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_12_LC_19_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41041),
            .lcout(M_this_scroll_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40329),
            .ce(N__27972),
            .sr(N__39763));
    defparam M_this_scroll_q_esr_15_LC_19_16_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_15_LC_19_16_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_15_LC_19_16_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_15_LC_19_16_0 (
            .in0(N__36458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_8_LC_19_16_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_8_LC_19_16_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_8_LC_19_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_8_LC_19_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35619),
            .lcout(M_this_scroll_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_9_LC_19_16_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_9_LC_19_16_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_9_LC_19_16_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_9_LC_19_16_2 (
            .in0(N__35512),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_11_LC_19_16_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_11_LC_19_16_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_11_LC_19_16_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_11_LC_19_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39506),
            .lcout(M_this_scroll_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_14_LC_19_16_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_14_LC_19_16_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_14_LC_19_16_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_14_LC_19_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36269),
            .lcout(M_this_scroll_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_13_LC_19_16_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_13_LC_19_16_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_13_LC_19_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_13_LC_19_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40599),
            .lcout(M_this_scroll_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam M_this_scroll_q_esr_10_LC_19_16_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_10_LC_19_16_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_10_LC_19_16_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_10_LC_19_16_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38784),
            .lcout(M_this_scroll_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40338),
            .ce(N__27973),
            .sr(N__39760));
    defparam \this_ppu.un1_M_hoffset_d_cry_0_c_LC_19_17_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_d_cry_0_c_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_d_cry_0_c_LC_19_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_d_cry_0_c_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(N__29345),
            .in2(N__29271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_19_17_0_),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_hoffset_q_esr_1_LC_19_17_1 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_1_LC_19_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_1_LC_19_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_1_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__27954),
            .in2(N__27910),
            .in3(N__27901),
            .lcout(\this_ppu.M_hoffset_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_0 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_1 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_2_LC_19_17_2 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_2_LC_19_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_2_LC_19_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_2_LC_19_17_2  (
            .in0(_gnd_net_),
            .in1(N__28379),
            .in2(N__28315),
            .in3(N__28306),
            .lcout(\this_ppu.M_hoffset_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_1 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_2 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_3_LC_19_17_3 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_3_LC_19_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_3_LC_19_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_3_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__28299),
            .in2(N__28225),
            .in3(N__28216),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_2 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_3 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_4_LC_19_17_4 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_4_LC_19_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_4_LC_19_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_4_LC_19_17_4  (
            .in0(_gnd_net_),
            .in1(N__28206),
            .in2(N__28159),
            .in3(N__28147),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_3 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_4 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_5_LC_19_17_5 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_5_LC_19_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_5_LC_19_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_5_LC_19_17_5  (
            .in0(_gnd_net_),
            .in1(N__28144),
            .in2(N__28131),
            .in3(N__28096),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_4 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_5 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_6_LC_19_17_6 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_6_LC_19_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_6_LC_19_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_6_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__28093),
            .in2(N__28086),
            .in3(N__28039),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_5 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_6 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_7_LC_19_17_7 .C_ON=1'b1;
    defparam \this_ppu.M_hoffset_q_esr_7_LC_19_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_7_LC_19_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_hoffset_q_esr_7_LC_19_17_7  (
            .in0(_gnd_net_),
            .in1(N__28036),
            .in2(N__28015),
            .in3(N__28006),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_d_cry_6 ),
            .carryout(\this_ppu.un1_M_hoffset_d_cry_7 ),
            .clk(N__40348),
            .ce(N__32058),
            .sr(N__39758));
    defparam \this_ppu.M_hoffset_q_esr_8_LC_19_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_hoffset_q_esr_8_LC_19_18_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_esr_8_LC_19_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.M_hoffset_q_esr_8_LC_19_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28003),
            .lcout(\this_ppu.M_hoffset_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40362),
            .ce(N__32050),
            .sr(N__39761));
    defparam \this_ppu.oam_cache.read_data_1_LC_19_20_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_1_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_1_LC_19_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_1_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40383),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_RNIPAFC_1_LC_19_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_RNIPAFC_1_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamidx_q_RNIPAFC_1_LC_19_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_oamidx_q_RNIPAFC_1_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(N__30300),
            .in2(_gnd_net_),
            .in3(N__28672),
            .lcout(),
            .ltout(\this_ppu.N_61_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_RNI8FTH1_0_LC_19_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_RNI8FTH1_0_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamidx_q_RNI8FTH1_0_LC_19_20_3 .LUT_INIT=16'b0000100000000100;
    LogicCell40 \this_ppu.M_oamidx_q_RNI8FTH1_0_LC_19_20_3  (
            .in0(N__29892),
            .in1(N__30037),
            .in2(N__28555),
            .in3(N__28740),
            .lcout(\this_ppu.N_769_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_3_LC_19_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_19_21_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_19_21_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_3_LC_19_21_2  (
            .in0(N__29847),
            .in1(N__33216),
            .in2(_gnd_net_),
            .in3(N__31548),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40394),
            .ce(),
            .sr(N__39768));
    defparam \this_ppu.M_state_q_2_LC_19_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_19_21_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_19_21_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.M_state_q_2_LC_19_21_5  (
            .in0(_gnd_net_),
            .in1(N__29521),
            .in2(_gnd_net_),
            .in3(N__29474),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40394),
            .ce(),
            .sr(N__39768));
    defparam \this_ppu.M_oamcurr_q_RNIMIF2_6_LC_19_22_1 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNIMIF2_6_LC_19_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNIMIF2_6_LC_19_22_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNIMIF2_6_LC_19_22_1  (
            .in0(N__28528),
            .in1(N__28462),
            .in2(N__28395),
            .in3(N__30163),
            .lcout(\this_ppu.N_779_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIUUIB7_6_LC_19_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIUUIB7_6_LC_19_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIUUIB7_6_LC_19_22_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_ppu.M_state_q_RNIUUIB7_6_LC_19_22_2  (
            .in0(N__29729),
            .in1(N__41398),
            .in2(N__28519),
            .in3(N__29827),
            .lcout(\this_ppu.un1_M_state_q_2_0 ),
            .ltout(\this_ppu.un1_M_state_q_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_2_LC_19_22_3 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_2_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_2_LC_19_22_3 .LUT_INIT=16'b1100011011001100;
    LogicCell40 \this_ppu.M_oamcurr_q_RNI6SKC7_2_LC_19_22_3  (
            .in0(N__28661),
            .in1(N__30070),
            .in2(N__28483),
            .in3(N__28728),
            .lcout(\this_ppu.M_oamcurr_q_RNI6SKC7Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_0_2_LC_19_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_0_2_LC_19_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNI6SKC7_0_2_LC_19_22_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNI6SKC7_0_2_LC_19_22_5  (
            .in0(N__28662),
            .in1(N__28729),
            .in2(N__30077),
            .in3(N__28617),
            .lcout(\this_ppu.un1_M_oamcurr_q_2_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_6_LC_19_22_7 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_6_LC_19_22_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamcurr_q_6_LC_19_22_7 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_oamcurr_q_6_LC_19_22_7  (
            .in0(N__28464),
            .in1(N__28438),
            .in2(N__28396),
            .in3(N__28408),
            .lcout(\this_ppu.M_oamcurr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40404),
            .ce(),
            .sr(N__28894));
    defparam \this_ppu.M_oamcurr_q_RNISRHKD_0_LC_19_23_1 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNISRHKD_0_LC_19_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNISRHKD_0_LC_19_23_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \this_ppu.M_oamcurr_q_RNISRHKD_0_LC_19_23_1  (
            .in0(N__28764),
            .in1(N__28734),
            .in2(_gnd_net_),
            .in3(N__28618),
            .lcout(\this_ppu.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI7KJ86_4_LC_19_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI7KJ86_4_LC_19_23_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI7KJ86_4_LC_19_23_2 .LUT_INIT=16'b0000100000001011;
    LogicCell40 \this_ppu.M_state_q_RNI7KJ86_4_LC_19_23_2  (
            .in0(N__29675),
            .in1(N__29415),
            .in2(N__39919),
            .in3(N__29998),
            .lcout(\this_ppu.N_329_0 ),
            .ltout(\this_ppu.N_329_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_RNIDG8LD_2_LC_19_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNIDG8LD_2_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNIDG8LD_2_LC_19_23_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNIDG8LD_2_LC_19_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28843),
            .in3(N__28839),
            .lcout(\this_ppu.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_RNI7SJLD_3_LC_19_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNI7SJLD_3_LC_19_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNI7SJLD_3_LC_19_23_4 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNI7SJLD_3_LC_19_23_4  (
            .in0(N__30178),
            .in1(N__28763),
            .in2(_gnd_net_),
            .in3(N__28805),
            .lcout(\this_ppu.N_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamcurr_q_RNIK5TKD_1_LC_19_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_oamcurr_q_RNIK5TKD_1_LC_19_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamcurr_q_RNIK5TKD_1_LC_19_23_5 .LUT_INIT=16'b1010000000101000;
    LogicCell40 \this_ppu.M_oamcurr_q_RNIK5TKD_1_LC_19_23_5  (
            .in0(N__28765),
            .in1(N__28733),
            .in2(N__28673),
            .in3(N__28619),
            .lcout(\this_ppu.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_19_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_19_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIPG425_1_LC_19_23_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIPG425_1_LC_19_23_6  (
            .in0(N__31799),
            .in1(N__31884),
            .in2(_gnd_net_),
            .in3(N__29999),
            .lcout(\this_ppu.un1_M_vaddress_q_c2 ),
            .ltout(\this_ppu.un1_M_vaddress_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_19_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_19_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_19_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_vaddress_q_RNIGPJH5_4_LC_19_23_7  (
            .in0(N__31716),
            .in1(N__31669),
            .in2(N__28579),
            .in3(N__31758),
            .lcout(\this_ppu.un1_M_vaddress_q_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_2_LC_19_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_2_LC_19_24_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamidx_q_2_LC_19_24_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \this_ppu.M_oamidx_q_2_LC_19_24_4  (
            .in0(N__30219),
            .in1(N__39911),
            .in2(N__30244),
            .in3(N__30021),
            .lcout(\this_ppu.M_oamidx_qZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40421),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_8_LC_19_24_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_8_LC_19_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_8_LC_19_24_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_8_LC_19_24_7  (
            .in0(N__28576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39328),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_9_LC_19_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_9_LC_19_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_9_LC_19_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_9_LC_19_25_0  (
            .in0(_gnd_net_),
            .in1(N__29083),
            .in2(_gnd_net_),
            .in3(N__39329),
            .lcout(M_this_oam_ram_write_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_14_LC_19_26_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_19_26_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_19_26_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_19_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36293),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40437),
            .ce(N__29064),
            .sr(N__39787));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_14_LC_19_28_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_14_LC_19_28_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_14_LC_19_28_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_14_LC_19_28_5  (
            .in0(_gnd_net_),
            .in1(N__29005),
            .in2(_gnd_net_),
            .in3(N__39368),
            .lcout(M_this_oam_ram_write_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_6_LC_20_12_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_6_LC_20_12_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_6_LC_20_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_6_LC_20_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28981),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40318),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_3_LC_20_14_3 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_3_LC_20_14_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_3_LC_20_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un20_i_a4_0_a3_0_a2_1_3_LC_20_14_3  (
            .in0(N__30359),
            .in1(N__36721),
            .in2(N__36797),
            .in3(N__30502),
            .lcout(),
            .ltout(\this_ppu.un20_i_a4_0_a3_0_a2_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_LC_20_14_4 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_LC_20_14_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \this_ppu.un20_i_a4_0_a3_0_a2_3_LC_20_14_4  (
            .in0(N__36667),
            .in1(_gnd_net_),
            .in2(N__28960),
            .in3(N__28956),
            .lcout(dma_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_12_LC_20_14_5.C_ON=1'b0;
    defparam M_this_state_q_12_LC_20_14_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_20_14_5.LUT_INIT=16'b0000000011001000;
    LogicCell40 M_this_state_q_12_LC_20_14_5 (
            .in0(N__40845),
            .in1(N__29254),
            .in2(N__30367),
            .in3(N__28906),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40330),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_i_LC_20_14_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_i_LC_20_14_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_i_LC_20_14_6 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_sn_m1_i_i_a3_i_i_LC_20_14_6  (
            .in0(N__36668),
            .in1(N__28957),
            .in2(_gnd_net_),
            .in3(N__40844),
            .lcout(N_260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_12_LC_20_14_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_12_LC_20_14_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_12_LC_20_14_7 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_a2_12_LC_20_14_7  (
            .in0(N__30360),
            .in1(N__32314),
            .in2(N__36798),
            .in3(N__30632),
            .lcout(\this_ppu.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_20_15_0.C_ON=1'b0;
    defparam M_this_state_q_11_LC_20_15_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_20_15_0.LUT_INIT=16'b1100100010001000;
    LogicCell40 M_this_state_q_11_LC_20_15_0 (
            .in0(N__36727),
            .in1(N__32121),
            .in2(N__30334),
            .in3(N__30501),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40339),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_12_LC_20_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_12_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_0_12_LC_20_15_2 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_0_12_LC_20_15_2  (
            .in0(N__39893),
            .in1(N__32193),
            .in2(_gnd_net_),
            .in3(N__36796),
            .lcout(\this_ppu.M_this_state_q_srsts_i_i_0_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_0_LC_20_15_5 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_0_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_3_0_LC_20_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un20_i_a4_0_a3_0_a2_3_0_LC_20_15_5  (
            .in0(N__30572),
            .in1(N__36726),
            .in2(N__36806),
            .in3(N__32262),
            .lcout(),
            .ltout(this_ppu_un20_i_a4_0_a3_0_a2_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI8K9F5_1_LC_20_15_6.C_ON=1'b0;
    defparam M_this_state_q_RNI8K9F5_1_LC_20_15_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI8K9F5_1_LC_20_15_6.LUT_INIT=16'b1000000011001100;
    LogicCell40 M_this_state_q_RNI8K9F5_1_LC_20_15_6 (
            .in0(N__30655),
            .in1(N__29248),
            .in2(N__29242),
            .in3(N__30508),
            .lcout(dma_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_11_LC_20_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_11_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_o2_11_LC_20_15_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_o2_11_LC_20_15_7  (
            .in0(_gnd_net_),
            .in1(N__40820),
            .in2(_gnd_net_),
            .in3(N__39892),
            .lcout(\this_ppu.N_328_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_10_LC_20_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_10_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_10_LC_20_16_0 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_1_10_LC_20_16_0  (
            .in0(N__40843),
            .in1(N__30499),
            .in2(N__32189),
            .in3(N__39904),
            .lcout(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_10_LC_20_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_10_LC_20_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_10_LC_20_16_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_10_LC_20_16_2  (
            .in0(_gnd_net_),
            .in1(N__30576),
            .in2(_gnd_net_),
            .in3(N__36731),
            .lcout(),
            .ltout(\this_ppu.N_414_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_20_16_3.C_ON=1'b0;
    defparam M_this_state_q_10_LC_20_16_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_20_16_3.LUT_INIT=16'b0000110010001100;
    LogicCell40 M_this_state_q_10_LC_20_16_3 (
            .in0(N__30500),
            .in1(N__29158),
            .in2(N__29152),
            .in3(N__30633),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40349),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_1_LC_20_16_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_ppu.M_state_q_RNO_0_1_LC_20_16_4  (
            .in0(N__41548),
            .in1(N__33223),
            .in2(N__29149),
            .in3(N__31549),
            .lcout(\this_ppu.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_20_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_20_17_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \this_ppu.M_state_q_1_LC_20_17_4  (
            .in0(N__29851),
            .in1(N__29362),
            .in2(N__41596),
            .in3(N__30019),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40363),
            .ce(),
            .sr(N__39757));
    defparam \this_ppu.M_hoffset_q_0_LC_20_18_5 .C_ON=1'b0;
    defparam \this_ppu.M_hoffset_q_0_LC_20_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_hoffset_q_0_LC_20_18_5 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \this_ppu.M_hoffset_q_0_LC_20_18_5  (
            .in0(N__29352),
            .in1(N__29820),
            .in2(N__29278),
            .in3(N__34135),
            .lcout(\this_ppu.hspr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40374),
            .ce(),
            .sr(N__39759));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_0_c_LC_20_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_0_c_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_0_c_LC_20_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_0_c_LC_20_19_0  (
            .in0(_gnd_net_),
            .in1(N__35785),
            .in2(N__34144),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_19_0_),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_LC_20_19_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_LC_20_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(N__35885),
            .in2(N__32653),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_0 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_LC_20_19_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_LC_20_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_LC_20_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(N__35325),
            .in2(N__34225),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_1 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_3_c_LC_20_19_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_3_c_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_3_c_LC_20_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_3_c_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(N__35020),
            .in2(N__33049),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_2 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_LC_20_19_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_LC_20_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_LC_20_19_4  (
            .in0(_gnd_net_),
            .in1(N__32978),
            .in2(N__32665),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_3 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_LC_20_19_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_LC_20_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_LC_20_19_5  (
            .in0(_gnd_net_),
            .in1(N__35178),
            .in2(N__32641),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_4 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_6_c_LC_20_19_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_6_c_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_6_c_LC_20_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_6_c_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(N__32860),
            .in2(N__32915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_5 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_LC_20_19_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_LC_20_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_LC_20_19_7  (
            .in0(_gnd_net_),
            .in1(N__31102),
            .in2(N__34302),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_2_cry_6 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_LC_20_20_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_LC_20_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_LC_20_20_0  (
            .in0(_gnd_net_),
            .in1(N__32677),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_20_0_),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNIH75J4_LC_20_20_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNIH75J4_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNIH75J4_LC_20_20_1 .LUT_INIT=16'b1111001101010001;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNIH75J4_LC_20_20_1  (
            .in0(N__32689),
            .in1(N__31108),
            .in2(N__32797),
            .in3(N__29737),
            .lcout(\this_ppu.N_242_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIPRKS1_1_LC_20_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIPRKS1_1_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIPRKS1_1_LC_20_20_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_ppu.M_state_q_RNIPRKS1_1_LC_20_20_2  (
            .in0(N__29813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39895),
            .lcout(\this_ppu.N_756_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_4_LC_20_20_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_4_LC_20_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_4_LC_20_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_4_LC_20_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29707),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40395),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_2_6_LC_20_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_2_6_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_2_6_LC_20_20_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_2_6_LC_20_20_4  (
            .in0(N__36973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37064),
            .lcout(\this_ppu.N_511 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIDM8L1_1_LC_20_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIDM8L1_1_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIDM8L1_1_LC_20_20_7 .LUT_INIT=16'b0000001011110010;
    LogicCell40 \this_ppu.M_state_q_RNIDM8L1_1_LC_20_20_7  (
            .in0(N__29514),
            .in1(N__29476),
            .in2(N__29436),
            .in3(N__29682),
            .lcout(\this_ppu.N_756_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNO_0_4_LC_20_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNO_0_4_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNO_0_4_LC_20_21_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_state_q_RNO_0_4_LC_20_21_4  (
            .in0(N__29518),
            .in1(N__29633),
            .in2(_gnd_net_),
            .in3(N__29581),
            .lcout(),
            .ltout(\this_ppu.N_799_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_20_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_20_21_5 .LUT_INIT=16'b0000110100000101;
    LogicCell40 \this_ppu.M_state_q_4_LC_20_21_5  (
            .in0(N__29530),
            .in1(N__29519),
            .in2(N__29479),
            .in3(N__29475),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40405),
            .ce(),
            .sr(N__39764));
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNI66L52_LC_20_21_6 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNI66L52_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNI66L52_LC_20_21_6 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_8_c_RNI66L52_LC_20_21_6  (
            .in0(N__29843),
            .in1(N__33215),
            .in2(_gnd_net_),
            .in3(N__31538),
            .lcout(\this_ppu.N_255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_voffset_q_0_LC_20_22_2 .C_ON=1'b0;
    defparam \this_ppu.M_voffset_q_0_LC_20_22_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_0_LC_20_22_2 .LUT_INIT=16'b0111101101001000;
    LogicCell40 \this_ppu.M_voffset_q_0_LC_20_22_2  (
            .in0(N__31880),
            .in1(N__29821),
            .in2(N__33187),
            .in3(N__34839),
            .lcout(\this_ppu.vspr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40415),
            .ce(),
            .sr(N__39769));
    defparam \this_ppu.M_vaddress_q_2_LC_20_23_2 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_2_LC_20_23_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_2_LC_20_23_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_2_LC_20_23_2  (
            .in0(N__31807),
            .in1(N__31768),
            .in2(N__31885),
            .in3(N__30025),
            .lcout(\this_ppu.M_vaddress_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.M_vaddress_q_3_LC_20_23_3 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_3_LC_20_23_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_3_LC_20_23_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_vaddress_q_3_LC_20_23_3  (
            .in0(N__31766),
            .in1(N__31718),
            .in2(_gnd_net_),
            .in3(N__29796),
            .lcout(\this_ppu.M_vaddress_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.M_vaddress_q_4_LC_20_23_4 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_4_LC_20_23_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_4_LC_20_23_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_4_LC_20_23_4  (
            .in0(N__29797),
            .in1(N__31673),
            .in2(N__31727),
            .in3(N__31767),
            .lcout(\this_ppu.M_vaddress_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.M_vaddress_q_7_LC_20_23_5 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_7_LC_20_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_7_LC_20_23_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \this_ppu.M_vaddress_q_7_LC_20_23_5  (
            .in0(N__29788),
            .in1(N__32077),
            .in2(N__31632),
            .in3(N__31577),
            .lcout(\this_ppu.M_vaddress_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.M_vaddress_q_5_LC_20_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_5_LC_20_23_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_5_LC_20_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.M_vaddress_q_5_LC_20_23_6  (
            .in0(_gnd_net_),
            .in1(N__31621),
            .in2(_gnd_net_),
            .in3(N__29786),
            .lcout(\this_ppu.M_vaddress_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.M_vaddress_q_6_LC_20_23_7 .C_ON=1'b0;
    defparam \this_ppu.M_vaddress_q_6_LC_20_23_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_vaddress_q_6_LC_20_23_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \this_ppu.M_vaddress_q_6_LC_20_23_7  (
            .in0(N__29787),
            .in1(_gnd_net_),
            .in2(N__31631),
            .in3(N__31576),
            .lcout(\this_ppu.M_vaddress_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40422),
            .ce(),
            .sr(N__29776));
    defparam \this_ppu.un1_M_oamidx_q_cry_0_c_LC_20_24_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oamidx_q_cry_0_c_LC_20_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oamidx_q_cry_0_c_LC_20_24_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oamidx_q_cry_0_c_LC_20_24_0  (
            .in0(_gnd_net_),
            .in1(N__41437),
            .in2(N__29884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_24_0_),
            .carryout(\this_ppu.un1_M_oamidx_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oamidx_q_cry_0_THRU_LUT4_0_LC_20_24_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oamidx_q_cry_0_THRU_LUT4_0_LC_20_24_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oamidx_q_cry_0_THRU_LUT4_0_LC_20_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oamidx_q_cry_0_THRU_LUT4_0_LC_20_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30299),
            .in3(N__30247),
            .lcout(\this_ppu.un1_M_oamidx_q_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oamidx_q_cry_0 ),
            .carryout(\this_ppu.un1_M_oamidx_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oamidx_q_cry_1_THRU_LUT4_0_LC_20_24_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oamidx_q_cry_1_THRU_LUT4_0_LC_20_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oamidx_q_cry_1_THRU_LUT4_0_LC_20_24_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oamidx_q_cry_1_THRU_LUT4_0_LC_20_24_2  (
            .in0(_gnd_net_),
            .in1(N__30218),
            .in2(_gnd_net_),
            .in3(N__30235),
            .lcout(\this_ppu.un1_M_oamidx_q_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oamidx_q_cry_1 ),
            .carryout(\this_ppu.un1_M_oamidx_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_3_LC_20_24_3 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_3_LC_20_24_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamidx_q_3_LC_20_24_3 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_ppu.M_oamidx_q_3_LC_20_24_3  (
            .in0(N__30024),
            .in1(N__39909),
            .in2(N__30120),
            .in3(N__30232),
            .lcout(\this_ppu.M_oamidx_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40429),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_RNIORUO_3_LC_20_24_5 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_RNIORUO_3_LC_20_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oamidx_q_RNIORUO_3_LC_20_24_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \this_ppu.M_oamidx_q_RNIORUO_3_LC_20_24_5  (
            .in0(N__30217),
            .in1(N__30182),
            .in2(N__30119),
            .in3(N__30081),
            .lcout(\this_ppu.M_state_q_srsts_0_a3_0_o2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oamidx_q_0_LC_20_24_6 .C_ON=1'b0;
    defparam \this_ppu.M_oamidx_q_0_LC_20_24_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oamidx_q_0_LC_20_24_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \this_ppu.M_oamidx_q_0_LC_20_24_6  (
            .in0(N__39910),
            .in1(N__41438),
            .in2(N__29885),
            .in3(N__30023),
            .lcout(\this_ppu.M_oamidx_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40429),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_2_LC_20_25_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_20_25_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_20_25_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_20_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38779),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40438),
            .ce(N__36015),
            .sr(N__39779));
    defparam M_this_data_tmp_q_esr_5_LC_20_25_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_20_25_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_20_25_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_20_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40607),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40438),
            .ce(N__36015),
            .sr(N__39779));
    defparam M_this_data_tmp_q_esr_19_LC_20_26_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_20_26_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_20_26_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_20_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39497),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40445),
            .ce(N__32437),
            .sr(N__39782));
    defparam M_this_data_tmp_q_esr_23_LC_20_26_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_20_26_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_20_26_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_20_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36487),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40445),
            .ce(N__32437),
            .sr(N__39782));
    defparam M_this_data_tmp_q_esr_17_LC_20_27_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_20_27_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_20_27_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_20_27_0 (
            .in0(N__35469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40450),
            .ce(N__32442),
            .sr(N__39788));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_7_LC_21_14_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_7_LC_21_14_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_7_LC_21_14_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_1_7_LC_21_14_0  (
            .in0(N__32266),
            .in1(N__30373),
            .in2(N__32194),
            .in3(N__39908),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_21_14_1.C_ON=1'b0;
    defparam M_this_state_q_7_LC_21_14_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_21_14_1.LUT_INIT=16'b1111000011100000;
    LogicCell40 M_this_state_q_7_LC_21_14_1 (
            .in0(N__30451),
            .in1(N__36670),
            .in2(N__30376),
            .in3(N__32267),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_7_LC_21_14_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_7_LC_21_14_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_7_LC_21_14_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_a2_1_7_LC_21_14_2  (
            .in0(N__36669),
            .in1(N__30539),
            .in2(_gnd_net_),
            .in3(N__30626),
            .lcout(\this_ppu.N_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a2_0_a2_0_2_LC_21_15_1 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a2_0_a2_0_2_LC_21_15_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a2_0_a2_0_2_LC_21_15_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.un20_i_a4_0_a2_0_a2_0_2_LC_21_15_1  (
            .in0(N__36775),
            .in1(N__30364),
            .in2(_gnd_net_),
            .in3(N__32260),
            .lcout(this_ppu_un20_i_a4_0_a2_0_a2_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_21_15_2.C_ON=1'b0;
    defparam M_this_state_q_4_LC_21_15_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_21_15_2.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_4_LC_21_15_2 (
            .in0(N__33790),
            .in1(N__32111),
            .in2(N__32346),
            .in3(N__30543),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40350),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_qlde_0_i_o2_0_LC_21_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_qlde_0_i_o2_0_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_qlde_0_i_o2_0_LC_21_15_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.M_this_data_count_qlde_0_i_o2_0_LC_21_15_3  (
            .in0(N__30366),
            .in1(N__32261),
            .in2(_gnd_net_),
            .in3(N__30498),
            .lcout(\this_ppu.N_341_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_13_LC_21_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_13_LC_21_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_i_0_1_13_LC_21_15_6 .LUT_INIT=16'b0000101100001010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_i_0_1_13_LC_21_15_6  (
            .in0(N__30365),
            .in1(N__40847),
            .in2(N__39921),
            .in3(N__36776),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_i_i_0_1Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_13_LC_21_15_7.C_ON=1'b0;
    defparam M_this_state_q_13_LC_21_15_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_21_15_7.LUT_INIT=16'b1111000010100000;
    LogicCell40 M_this_state_q_13_LC_21_15_7 (
            .in0(N__36777),
            .in1(_gnd_net_),
            .in2(N__30337),
            .in3(N__30330),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40350),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_5_LC_21_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_5_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_5_LC_21_16_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_5_LC_21_16_0  (
            .in0(N__30571),
            .in1(_gnd_net_),
            .in2(N__32122),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_ppu.N_424_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_21_16_1.C_ON=1'b0;
    defparam M_this_state_q_5_LC_21_16_1.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_21_16_1.LUT_INIT=16'b1111100011110000;
    LogicCell40 M_this_state_q_5_LC_21_16_1 (
            .in0(N__36985),
            .in1(N__37078),
            .in2(N__30667),
            .in3(N__33789),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40364),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_data_count_qlde_0_i_a2_LC_21_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_data_count_qlde_0_i_a2_LC_21_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_data_count_qlde_0_i_a2_LC_21_16_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \this_ppu.M_this_data_count_qlde_0_i_a2_LC_21_16_2  (
            .in0(N__30645),
            .in1(N__32185),
            .in2(_gnd_net_),
            .in3(N__30627),
            .lcout(\this_ppu.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI1G0L_1_LC_21_16_3.C_ON=1'b0;
    defparam M_this_state_q_RNI1G0L_1_LC_21_16_3.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI1G0L_1_LC_21_16_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 M_this_state_q_RNI1G0L_1_LC_21_16_3 (
            .in0(N__36508),
            .in1(N__36683),
            .in2(_gnd_net_),
            .in3(N__32626),
            .lcout(M_this_state_q_RNI1G0LZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_1_0_0_LC_21_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_1_0_0_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_1_0_0_LC_21_16_4 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_i_1_0_0_LC_21_16_4  (
            .in0(N__32107),
            .in1(N__32563),
            .in2(N__30649),
            .in3(N__30628),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_i_1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a2_0_o2_2_LC_21_16_5 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a2_0_o2_2_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a2_0_o2_2_LC_21_16_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_ppu.un20_i_a4_0_a2_0_o2_2_LC_21_16_5  (
            .in0(N__32301),
            .in1(N__30570),
            .in2(_gnd_net_),
            .in3(N__30538),
            .lcout(N_311_0),
            .ltout(N_311_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNI244K2_10_LC_21_16_6.C_ON=1'b0;
    defparam M_this_state_q_RNI244K2_10_LC_21_16_6.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNI244K2_10_LC_21_16_6.LUT_INIT=16'b0001010100111111;
    LogicCell40 M_this_state_q_RNI244K2_10_LC_21_16_6 (
            .in0(N__32227),
            .in1(N__30517),
            .in2(N__30511),
            .in3(N__30466),
            .lcout(M_this_state_q_RNI244K2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIR71E_10_LC_21_16_7.C_ON=1'b0;
    defparam M_this_state_q_RNIR71E_10_LC_21_16_7.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIR71E_10_LC_21_16_7.LUT_INIT=16'b0000000000110011;
    LogicCell40 M_this_state_q_RNIR71E_10_LC_21_16_7 (
            .in0(_gnd_net_),
            .in1(N__36722),
            .in2(_gnd_net_),
            .in3(N__30494),
            .lcout(M_this_state_q_RNIR71EZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.hspr_cry_0_c_inv_LC_21_17_0 .C_ON=1'b1;
    defparam \this_ppu.hspr_cry_0_c_inv_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.hspr_cry_0_c_inv_LC_21_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.hspr_cry_0_c_inv_LC_21_17_0  (
            .in0(N__35784),
            .in1(N__34134),
            .in2(N__30460),
            .in3(_gnd_net_),
            .lcout(\this_ppu.hspr_cry_0_c_inv_RNI1203 ),
            .ltout(),
            .carryin(bfn_21_17_0_),
            .carryout(\this_ppu.hspr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.hspr_cry_0_c_RNISEIH1_LC_21_17_1 .C_ON=1'b1;
    defparam \this_ppu.hspr_cry_0_c_RNISEIH1_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.hspr_cry_0_c_RNISEIH1_LC_21_17_1 .LUT_INIT=16'b1100100110011100;
    LogicCell40 \this_ppu.hspr_cry_0_c_RNISEIH1_LC_21_17_1  (
            .in0(N__34966),
            .in1(N__35886),
            .in2(N__30676),
            .in3(N__30895),
            .lcout(M_this_ppu_spr_addr_1),
            .ltout(),
            .carryin(\this_ppu.hspr_cry_0 ),
            .carryout(\this_ppu.hspr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.hspr_cry_1_c_RNI6K8I1_LC_21_17_2 .C_ON=1'b0;
    defparam \this_ppu.hspr_cry_1_c_RNI6K8I1_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.hspr_cry_1_c_RNI6K8I1_LC_21_17_2 .LUT_INIT=16'b1001110011001001;
    LogicCell40 \this_ppu.hspr_cry_1_c_RNI6K8I1_LC_21_17_2  (
            .in0(N__34967),
            .in1(N__35324),
            .in2(N__36586),
            .in3(N__30892),
            .lcout(M_this_ppu_spr_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_21_17_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_21_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_21_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIUU07_9_LC_21_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35848),
            .lcout(\this_ppu.M_oam_cache_read_data_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_inv_LC_21_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_inv_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_inv_LC_21_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_0_c_inv_LC_21_18_0  (
            .in0(_gnd_net_),
            .in1(N__35782),
            .in2(N__32538),
            .in3(N__34124),
            .lcout(\this_ppu.M_hoffset_q_i_0 ),
            .ltout(),
            .carryin(bfn_21_18_0_),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_inv_LC_21_18_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_inv_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_inv_LC_21_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_1_c_inv_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__35846),
            .in2(N__32520),
            .in3(N__35887),
            .lcout(\this_ppu.M_hoffset_q_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_0 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_inv_LC_21_18_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_inv_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_inv_LC_21_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_2_c_inv_LC_21_18_2  (
            .in0(_gnd_net_),
            .in1(N__36582),
            .in2(N__32502),
            .in3(N__35332),
            .lcout(\this_ppu.M_hoffset_q_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_1 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_inv_LC_21_18_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_inv_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_inv_LC_21_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_3_c_inv_LC_21_18_3  (
            .in0(_gnd_net_),
            .in1(N__35931),
            .in2(N__32481),
            .in3(N__33050),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_0 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_2 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_inv_LC_21_18_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_inv_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_inv_LC_21_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_4_c_inv_LC_21_18_4  (
            .in0(_gnd_net_),
            .in1(N__35077),
            .in2(N__32463),
            .in3(N__32985),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_3 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_inv_LC_21_18_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_inv_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_inv_LC_21_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_5_c_inv_LC_21_18_5  (
            .in0(_gnd_net_),
            .in1(N__35124),
            .in2(N__32739),
            .in3(N__35174),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_4 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_inv_LC_21_18_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_inv_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_inv_LC_21_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_6_c_inv_LC_21_18_6  (
            .in0(_gnd_net_),
            .in1(N__34427),
            .in2(N__32721),
            .in3(N__32902),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_5 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_inv_LC_21_18_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_inv_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_inv_LC_21_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_7_c_inv_LC_21_18_7  (
            .in0(_gnd_net_),
            .in1(N__32703),
            .in2(N__34368),
            .in3(N__34286),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_2_cry_6 ),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_inv_LC_21_19_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_inv_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_inv_LC_21_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_2_cry_8_c_inv_LC_21_19_0  (
            .in0(_gnd_net_),
            .in1(N__31117),
            .in2(_gnd_net_),
            .in3(N__32822),
            .lcout(\this_ppu.M_hoffset_q_i_8 ),
            .ltout(),
            .carryin(bfn_21_19_0_),
            .carryout(\this_ppu.un1_M_hoffset_q_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_RNITUI32_LC_21_19_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_RNITUI32_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_2_cry_8_c_RNITUI32_LC_21_19_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_2_cry_8_c_RNITUI32_LC_21_19_1  (
            .in0(N__34367),
            .in1(N__34393),
            .in2(_gnd_net_),
            .in3(N__31111),
            .lcout(\this_ppu.vspr12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNO_LC_21_19_3 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNO_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNO_LC_21_19_3 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNO_LC_21_19_3  (
            .in0(N__34366),
            .in1(N__34392),
            .in2(_gnd_net_),
            .in3(N__34296),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_2_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_0_c_LC_21_20_0 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_LC_21_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_0_c_LC_21_20_0  (
            .in0(_gnd_net_),
            .in1(N__39061),
            .in2(N__34857),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_20_0_),
            .carryout(\this_ppu.un1_oam_data_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_1_c_LC_21_20_1 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_LC_21_20_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_1_c_LC_21_20_1  (
            .in0(_gnd_net_),
            .in1(N__39010),
            .in2(N__33106),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_0 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_2_c_LC_21_20_2 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_LC_21_20_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_2_c_LC_21_20_2  (
            .in0(_gnd_net_),
            .in1(N__38389),
            .in2(N__33538),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_1 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_3_c_LC_21_20_3 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_LC_21_20_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_3_c_LC_21_20_3  (
            .in0(_gnd_net_),
            .in1(N__38182),
            .in2(N__33489),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_2 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_4_c_LC_21_20_4 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_LC_21_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_LC_21_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_4_c_LC_21_20_4  (
            .in0(_gnd_net_),
            .in1(N__38596),
            .in2(N__33438),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_3 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_5_c_LC_21_20_5 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_LC_21_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_5_c_LC_21_20_5  (
            .in0(_gnd_net_),
            .in1(N__32746),
            .in2(N__33390),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_4 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_6_c_LC_21_20_6 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_LC_21_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_6_c_LC_21_20_6  (
            .in0(_gnd_net_),
            .in1(N__32764),
            .in2(N__33345),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_5 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_7_c_LC_21_20_7 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_7_c_LC_21_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_7_c_LC_21_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_7_c_LC_21_20_7  (
            .in0(_gnd_net_),
            .in1(N__32752),
            .in2(N__33291),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_6 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_8_c_LC_21_21_0 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_LC_21_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_8_c_LC_21_21_0  (
            .in0(_gnd_net_),
            .in1(N__32758),
            .in2(N__33250),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_21_0_),
            .carryout(\this_ppu.un1_oam_data_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_8_THRU_LUT4_0_LC_21_21_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_8_THRU_LUT4_0_LC_21_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_8_THRU_LUT4_0_LC_21_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_8_THRU_LUT4_0_LC_21_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31552),
            .lcout(\this_ppu.un1_oam_data_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vspr_cry_0_c_inv_LC_21_22_0 .C_ON=1'b1;
    defparam \this_ppu.vspr_cry_0_c_inv_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vspr_cry_0_c_inv_LC_21_22_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.vspr_cry_0_c_inv_LC_21_22_0  (
            .in0(_gnd_net_),
            .in1(N__34843),
            .in2(N__31522),
            .in3(N__35401),
            .lcout(\this_ppu.vspr_cry_0_c_inv_RNIFK43 ),
            .ltout(),
            .carryin(bfn_21_22_0_),
            .carryout(\this_ppu.vspr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vspr_cry_0_c_RNI75JG1_LC_21_22_1 .C_ON=1'b1;
    defparam \this_ppu.vspr_cry_0_c_RNI75JG1_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vspr_cry_0_c_RNI75JG1_LC_21_22_1 .LUT_INIT=16'b1100100110011100;
    LogicCell40 \this_ppu.vspr_cry_0_c_RNI75JG1_LC_21_22_1  (
            .in0(N__34940),
            .in1(N__33102),
            .in2(N__31912),
            .in3(N__31315),
            .lcout(M_this_ppu_spr_addr_4),
            .ltout(),
            .carryin(\this_ppu.vspr_cry_0 ),
            .carryout(\this_ppu.vspr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.vspr_cry_1_c_RNIA9KG1_LC_21_22_2 .C_ON=1'b0;
    defparam \this_ppu.vspr_cry_1_c_RNIA9KG1_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.vspr_cry_1_c_RNIA9KG1_LC_21_22_2 .LUT_INIT=16'b1101001011100001;
    LogicCell40 \this_ppu.vspr_cry_1_c_RNIA9KG1_LC_21_22_2  (
            .in0(N__32770),
            .in1(N__34941),
            .in2(N__33537),
            .in3(N__31312),
            .lcout(M_this_ppu_spr_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_21_22_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_21_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNID8M7_17_LC_21_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31891),
            .lcout(\this_ppu.M_oam_cache_read_data_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_17_LC_21_22_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_17_LC_21_22_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_17_LC_21_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_17_LC_21_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31903),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40423),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_d_cry_0_c_LC_21_23_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_d_cry_0_c_LC_21_23_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_d_cry_0_c_LC_21_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_voffset_d_cry_0_c_LC_21_23_0  (
            .in0(_gnd_net_),
            .in1(N__31876),
            .in2(N__33180),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_23_0_),
            .carryout(\this_ppu.un1_M_voffset_d_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_voffset_q_esr_1_LC_21_23_1 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_1_LC_21_23_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_1_LC_21_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_1_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(N__31806),
            .in2(N__33163),
            .in3(N__31771),
            .lcout(\this_ppu.M_voffset_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_0 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_1 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_2_LC_21_23_2 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_2_LC_21_23_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_2_LC_21_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_2_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(N__31757),
            .in2(N__33655),
            .in3(N__31741),
            .lcout(\this_ppu.M_voffset_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_1 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_2 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_3_LC_21_23_3 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_3_LC_21_23_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_3_LC_21_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_3_LC_21_23_3  (
            .in0(_gnd_net_),
            .in1(N__31717),
            .in2(N__33145),
            .in3(N__31690),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_2 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_3 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_4_LC_21_23_4 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_4_LC_21_23_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_4_LC_21_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_4_LC_21_23_4  (
            .in0(_gnd_net_),
            .in1(N__33136),
            .in2(N__31677),
            .in3(N__31645),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_3 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_4 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_5_LC_21_23_5 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_5_LC_21_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_5_LC_21_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_5_LC_21_23_5  (
            .in0(_gnd_net_),
            .in1(N__31617),
            .in2(N__33154),
            .in3(N__31597),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_4 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_5 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_6_LC_21_23_6 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_6_LC_21_23_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_6_LC_21_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_6_LC_21_23_6  (
            .in0(_gnd_net_),
            .in1(N__33130),
            .in2(N__31581),
            .in3(N__32080),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_5 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_6 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_7_LC_21_23_7 .C_ON=1'b1;
    defparam \this_ppu.M_voffset_q_esr_7_LC_21_23_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_7_LC_21_23_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_voffset_q_esr_7_LC_21_23_7  (
            .in0(_gnd_net_),
            .in1(N__32076),
            .in2(N__33124),
            .in3(N__32065),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_d_cry_6 ),
            .carryout(\this_ppu.un1_M_voffset_d_cry_7 ),
            .clk(N__40430),
            .ce(N__32057),
            .sr(N__39770));
    defparam \this_ppu.M_voffset_q_esr_8_LC_21_24_0 .C_ON=1'b0;
    defparam \this_ppu.M_voffset_q_esr_8_LC_21_24_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_voffset_q_esr_8_LC_21_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.M_voffset_q_esr_8_LC_21_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32062),
            .lcout(\this_ppu.M_voffset_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40439),
            .ce(N__32059),
            .sr(N__39773));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_2_LC_21_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_2_LC_21_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_2_LC_21_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_2_LC_21_25_0  (
            .in0(N__39348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32011),
            .lcout(M_this_oam_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_16_LC_21_25_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_16_LC_21_25_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_16_LC_21_25_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_16_LC_21_25_4  (
            .in0(N__39347),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31993),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_5_LC_21_25_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_5_LC_21_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_5_LC_21_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_5_LC_21_25_5  (
            .in0(_gnd_net_),
            .in1(N__31966),
            .in2(_gnd_net_),
            .in3(N__39349),
            .lcout(M_this_oam_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_15_LC_21_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_15_LC_21_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_15_LC_21_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_15_LC_21_25_7  (
            .in0(_gnd_net_),
            .in1(N__31948),
            .in2(_gnd_net_),
            .in3(N__39346),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_19_LC_21_26_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_19_LC_21_26_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_19_LC_21_26_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_19_LC_21_26_0  (
            .in0(N__39372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31930),
            .lcout(M_this_oam_ram_write_data_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_0_LC_21_27_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_21_27_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_21_27_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_21_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35563),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40454),
            .ce(N__36028),
            .sr(N__39783));
    defparam M_this_data_tmp_q_esr_22_LC_21_28_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_21_28_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_21_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_21_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36307),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40460),
            .ce(N__32446),
            .sr(N__39789));
    defparam \this_spr_ram.mem_radreg_13_LC_22_11_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_13_LC_22_11_0 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_13_LC_22_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_13_LC_22_11_0  (
            .in0(N__34171),
            .in1(N__32365),
            .in2(_gnd_net_),
            .in3(N__34981),
            .lcout(\this_spr_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40323),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_i_1_6_LC_22_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_i_1_6_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_i_1_6_LC_22_15_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_i_1_6_LC_22_15_2  (
            .in0(N__39902),
            .in1(N__33751),
            .in2(N__32350),
            .in3(N__36885),
            .lcout(),
            .ltout(\this_ppu.M_this_state_q_srsts_0_i_0_i_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_22_15_3.C_ON=1'b0;
    defparam M_this_state_q_6_LC_22_15_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_22_15_3.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_6_LC_22_15_3 (
            .in0(N__33715),
            .in1(N__32123),
            .in2(N__32317),
            .in3(N__32309),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40365),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_LC_22_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_LC_22_15_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_LC_22_15_7 .LUT_INIT=16'b0000000010100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_0_a2_1_LC_22_15_7  (
            .in0(N__36519),
            .in1(N__40846),
            .in2(N__36893),
            .in3(N__39901),
            .lcout(\this_ppu.N_416 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_22_16_0.C_ON=1'b0;
    defparam M_this_state_q_2_LC_22_16_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_22_16_0.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_2_LC_22_16_0 (
            .in0(N__32132),
            .in1(N__33778),
            .in2(N__32601),
            .in3(N__33802),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40375),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_1_LC_22_16_2 .C_ON=1'b0;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_1_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un20_i_a4_0_a3_0_a2_1_1_LC_22_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un20_i_a4_0_a3_0_a2_1_1_LC_22_16_2  (
            .in0(N__32302),
            .in1(N__32586),
            .in2(N__32629),
            .in3(N__32268),
            .lcout(this_ppu_un20_i_a4_0_a3_0_a2_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_3_6_LC_22_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_3_6_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_3_6_LC_22_16_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_3_6_LC_22_16_5  (
            .in0(N__41269),
            .in1(N__32221),
            .in2(_gnd_net_),
            .in3(N__32184),
            .lcout(\this_ppu.N_916 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_22_16_6.C_ON=1'b0;
    defparam M_this_state_q_3_LC_22_16_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_22_16_6.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_3_LC_22_16_6 (
            .in0(N__32625),
            .in1(N__33796),
            .in2(N__32137),
            .in3(N__33779),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40375),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIKV6G1_2_LC_22_17_0.C_ON=1'b0;
    defparam M_this_state_q_RNIKV6G1_2_LC_22_17_0.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIKV6G1_2_LC_22_17_0.LUT_INIT=16'b1010111010101010;
    LogicCell40 M_this_state_q_RNIKV6G1_2_LC_22_17_0 (
            .in0(N__39884),
            .in1(N__32628),
            .in2(N__32597),
            .in3(N__40848),
            .lcout(N_1318_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_a2_1_0_LC_22_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_a2_1_0_LC_22_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_i_a2_1_0_LC_22_17_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_i_a2_1_0_LC_22_17_5  (
            .in0(N__32627),
            .in1(N__32590),
            .in2(N__36518),
            .in3(N__39885),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0 ),
            .ltout(\this_ppu.M_this_state_q_srsts_0_i_i_a2_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_22_17_6.C_ON=1'b0;
    defparam M_this_state_q_0_LC_22_17_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_22_17_6.LUT_INIT=16'b1111111101001100;
    LogicCell40 M_this_state_q_0_LC_22_17_6 (
            .in0(N__36843),
            .in1(N__36886),
            .in2(N__32557),
            .in3(N__32554),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40384),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_22_17_7.C_ON=1'b0;
    defparam M_this_state_q_1_LC_22_17_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_22_17_7.LUT_INIT=16'b1100110111001100;
    LogicCell40 M_this_state_q_1_LC_22_17_7 (
            .in0(N__36966),
            .in1(N__32548),
            .in2(N__37077),
            .in3(N__33774),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40384),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_LC_22_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_LC_22_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_0_c_LC_22_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_0_c_LC_22_18_0  (
            .in0(_gnd_net_),
            .in1(N__35783),
            .in2(N__32539),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_18_0_),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_LC_22_18_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_1_c_LC_22_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_1_c_LC_22_18_1  (
            .in0(_gnd_net_),
            .in1(N__35847),
            .in2(N__32521),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_0 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_LC_22_18_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_2_c_LC_22_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_2_c_LC_22_18_2  (
            .in0(_gnd_net_),
            .in1(N__36581),
            .in2(N__32503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_1 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_LC_22_18_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_3_c_LC_22_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_3_c_LC_22_18_3  (
            .in0(_gnd_net_),
            .in1(N__35932),
            .in2(N__32485),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_2 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_LC_22_18_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_4_c_LC_22_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_4_c_LC_22_18_4  (
            .in0(_gnd_net_),
            .in1(N__35072),
            .in2(N__32464),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_3 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_LC_22_18_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_LC_22_18_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_5_c_LC_22_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_5_c_LC_22_18_5  (
            .in0(_gnd_net_),
            .in1(N__35125),
            .in2(N__32740),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_4 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_LC_22_18_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_LC_22_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_6_c_LC_22_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_6_c_LC_22_18_6  (
            .in0(_gnd_net_),
            .in1(N__34428),
            .in2(N__32722),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_5 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_LC_22_18_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_LC_22_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_7_c_LC_22_18_7  (
            .in0(_gnd_net_),
            .in1(N__32704),
            .in2(N__34369),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_hoffset_q_cry_6 ),
            .carryout(\this_ppu.un1_M_hoffset_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_RNIB1P42_LC_22_19_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_RNIB1P42_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_hoffset_q_cry_7_c_RNIB1P42_LC_22_19_0 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_ppu.un1_M_hoffset_q_cry_7_c_RNIB1P42_LC_22_19_0  (
            .in0(N__34386),
            .in1(N__34354),
            .in2(_gnd_net_),
            .in3(N__32692),
            .lcout(\this_ppu.vspr16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_RNO_LC_22_19_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_RNO_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_RNO_LC_22_19_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_8_c_RNO_LC_22_19_1  (
            .in0(_gnd_net_),
            .in1(N__34344),
            .in2(_gnd_net_),
            .in3(N__34385),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_ac0_13_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNO_LC_22_19_3 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNO_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNO_LC_22_19_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNO_LC_22_19_3  (
            .in0(N__32826),
            .in1(N__34343),
            .in2(_gnd_net_),
            .in3(N__34384),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNO_LC_22_19_4 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNO_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNO_LC_22_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNO_LC_22_19_4  (
            .in0(N__32989),
            .in1(N__35065),
            .in2(_gnd_net_),
            .in3(N__35229),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_2_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNO_LC_22_19_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNO_LC_22_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNO_LC_22_19_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNO_LC_22_19_6  (
            .in0(N__35898),
            .in1(N__35826),
            .in2(_gnd_net_),
            .in3(N__35761),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_2_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNO_LC_22_19_7 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNO_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNO_LC_22_19_7 .LUT_INIT=16'b1010000001011111;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNO_LC_22_19_7  (
            .in0(N__35230),
            .in1(N__35182),
            .in2(N__35073),
            .in3(N__35117),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_2_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNO_LC_22_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNO_LC_22_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNO_LC_22_20_0 .LUT_INIT=16'b1010000001011111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_6_c_RNO_LC_22_20_0  (
            .in0(N__35693),
            .in1(_gnd_net_),
            .in2(N__34499),
            .in3(N__34558),
            .lcout(\this_ppu.un1_oam_data_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNO_LC_22_20_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNO_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_8_c_RNO_LC_22_20_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_8_c_RNO_LC_22_20_1  (
            .in0(N__34560),
            .in1(N__34495),
            .in2(N__35680),
            .in3(N__35695),
            .lcout(\this_ppu.un1_oam_data_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_7_c_RNO_LC_22_20_2 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_7_c_RNO_LC_22_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_7_c_RNO_LC_22_20_2 .LUT_INIT=16'b1001001100110011;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_7_c_RNO_LC_22_20_2  (
            .in0(N__35694),
            .in1(N__35675),
            .in2(N__34500),
            .in3(N__34559),
            .lcout(\this_ppu.un1_oam_data_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_14_LC_22_20_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_14_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_14_LC_22_20_3 .LUT_INIT=16'b1000011100001111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI3DGK1_14_LC_22_20_3  (
            .in0(N__35228),
            .in1(N__35108),
            .in2(N__34429),
            .in3(N__35063),
            .lcout(\this_ppu.read_data_RNI3DGK1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNO_LC_22_20_5 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNO_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNO_LC_22_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_5_c_RNO_LC_22_20_5  (
            .in0(_gnd_net_),
            .in1(N__34488),
            .in2(_gnd_net_),
            .in3(N__35692),
            .lcout(\this_ppu.un1_oam_data_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNO_LC_22_20_7 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNO_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNO_LC_22_20_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNO_LC_22_20_7  (
            .in0(N__35227),
            .in1(N__32990),
            .in2(_gnd_net_),
            .in3(N__35062),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_0_c_LC_22_21_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_0_c_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_0_c_LC_22_21_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_0_c_LC_22_21_0  (
            .in0(_gnd_net_),
            .in1(N__35753),
            .in2(N__34154),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_21_0_),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_LC_22_21_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_LC_22_21_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_LC_22_21_1  (
            .in0(_gnd_net_),
            .in1(N__35897),
            .in2(N__35704),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_0 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_LC_22_21_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_LC_22_21_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_LC_22_21_2  (
            .in0(_gnd_net_),
            .in1(N__35333),
            .in2(N__35275),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_1 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_3_c_LC_22_21_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_3_c_LC_22_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_3_c_LC_22_21_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_3_c_LC_22_21_3  (
            .in0(_gnd_net_),
            .in1(N__35013),
            .in2(N__33063),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_2 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_LC_22_21_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_LC_22_21_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_4_c_LC_22_21_4  (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(N__32994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_3 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_LC_22_21_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_LC_22_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_LC_22_21_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_LC_22_21_5  (
            .in0(_gnd_net_),
            .in1(N__35026),
            .in2(N__35199),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_4 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_6_c_LC_22_21_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_6_c_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_6_c_LC_22_21_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_6_c_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__32919),
            .in2(N__32856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_5 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_LC_22_21_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_LC_22_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_LC_22_21_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_LC_22_21_7  (
            .in0(_gnd_net_),
            .in1(N__34300),
            .in2(N__34237),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_read_data_3_cry_6 ),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_LC_22_22_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_LC_22_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_8_c_LC_22_22_0  (
            .in0(_gnd_net_),
            .in1(N__32839),
            .in2(N__32830),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_22_22_0_),
            .carryout(\this_ppu.un1_M_oam_cache_read_data_3_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_LUT4_0_LC_22_22_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_LUT4_0_LC_22_22_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_LUT4_0_LC_22_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_LUT4_0_LC_22_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32800),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_18_LC_22_22_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_18_LC_22_22_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_18_LC_22_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_18_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32782),
            .lcout(\this_ppu.M_oam_cache_read_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40431),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_0_LC_22_23_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_0_LC_22_23_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_0_LC_22_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_0_LC_22_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35569),
            .lcout(M_this_scroll_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_1_LC_22_23_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_1_LC_22_23_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_1_LC_22_23_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_1_LC_22_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35475),
            .lcout(M_this_scroll_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_5_LC_22_23_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_5_LC_22_23_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_5_LC_22_23_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_5_LC_22_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40574),
            .lcout(M_this_scroll_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_3_LC_22_23_3.C_ON=1'b0;
    defparam M_this_scroll_q_esr_3_LC_22_23_3.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_3_LC_22_23_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_3_LC_22_23_3 (
            .in0(N__39454),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_4_LC_22_23_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_4_LC_22_23_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_4_LC_22_23_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_4_LC_22_23_4 (
            .in0(N__41016),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_6_LC_22_23_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_6_LC_22_23_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_6_LC_22_23_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_6_LC_22_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36262),
            .lcout(M_this_scroll_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam M_this_scroll_q_esr_7_LC_22_23_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_7_LC_22_23_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_7_LC_22_23_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 M_this_scroll_q_esr_7_LC_22_23_7 (
            .in0(_gnd_net_),
            .in1(N__36462),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40440),
            .ce(N__33633),
            .sr(N__39765));
    defparam \this_ppu.un1_M_voffset_q_cry_0_c_inv_LC_22_24_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_0_c_inv_LC_22_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_0_c_inv_LC_22_24_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_0_c_inv_LC_22_24_0  (
            .in0(_gnd_net_),
            .in1(N__39057),
            .in2(N__33115),
            .in3(N__34850),
            .lcout(\this_ppu.M_voffset_q_i_0 ),
            .ltout(),
            .carryin(bfn_22_24_0_),
            .carryout(\this_ppu.un1_M_voffset_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_1_c_inv_LC_22_24_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_1_c_inv_LC_22_24_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_1_c_inv_LC_22_24_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_1_c_inv_LC_22_24_1  (
            .in0(_gnd_net_),
            .in1(N__39103),
            .in2(N__33082),
            .in3(N__33098),
            .lcout(\this_ppu.M_voffset_q_i_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_0 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_2_c_inv_LC_22_24_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_2_c_inv_LC_22_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_2_c_inv_LC_22_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_2_c_inv_LC_22_24_2  (
            .in0(_gnd_net_),
            .in1(N__38441),
            .in2(N__33511),
            .in3(N__33527),
            .lcout(\this_ppu.M_voffset_q_i_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_1 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_3_c_inv_LC_22_24_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_3_c_inv_LC_22_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_3_c_inv_LC_22_24_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_3_c_inv_LC_22_24_3  (
            .in0(_gnd_net_),
            .in1(N__38565),
            .in2(N__33457),
            .in3(N__33476),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_2 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_4_c_inv_LC_22_24_4 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_4_c_inv_LC_22_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_4_c_inv_LC_22_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_4_c_inv_LC_22_24_4  (
            .in0(_gnd_net_),
            .in1(N__38508),
            .in2(N__33406),
            .in3(N__33425),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_3 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_5_c_inv_LC_22_24_5 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_5_c_inv_LC_22_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_5_c_inv_LC_22_24_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_5_c_inv_LC_22_24_5  (
            .in0(_gnd_net_),
            .in1(N__34484),
            .in2(N__33358),
            .in3(N__33377),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_7 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_4 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_6_c_inv_LC_22_24_6 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_6_c_inv_LC_22_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_6_c_inv_LC_22_24_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_6_c_inv_LC_22_24_6  (
            .in0(_gnd_net_),
            .in1(N__34554),
            .in2(N__33307),
            .in3(N__33326),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_8 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_5 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_7_c_inv_LC_22_24_7 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_7_c_inv_LC_22_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_7_c_inv_LC_22_24_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_7_c_inv_LC_22_24_7  (
            .in0(_gnd_net_),
            .in1(N__35671),
            .in2(N__33259),
            .in3(N__33278),
            .lcout(\this_ppu.M_this_ppu_map_addr_i_9 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_voffset_q_cry_6 ),
            .carryout(\this_ppu.un1_M_voffset_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_inv_LC_22_25_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_inv_LC_22_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_inv_LC_22_25_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_8_c_inv_LC_22_25_0  (
            .in0(_gnd_net_),
            .in1(N__33232),
            .in2(_gnd_net_),
            .in3(N__33243),
            .lcout(\this_ppu.M_voffset_q_i_8 ),
            .ltout(),
            .carryin(bfn_22_25_0_),
            .carryout(\this_ppu.un1_M_voffset_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_RNICN6N1_LC_22_25_1 .C_ON=1'b0;
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_RNICN6N1_LC_22_25_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_voffset_q_cry_8_c_RNICN6N1_LC_22_25_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_ppu.un1_M_voffset_q_cry_8_c_RNICN6N1_LC_22_25_1  (
            .in0(N__38209),
            .in1(N__38044),
            .in2(_gnd_net_),
            .in3(N__33226),
            .lcout(\this_ppu.M_state_d14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_24_LC_22_25_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_24_LC_22_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_24_LC_22_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_24_LC_22_25_2  (
            .in0(_gnd_net_),
            .in1(N__35598),
            .in2(_gnd_net_),
            .in3(N__39333),
            .lcout(N_433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_29_LC_22_25_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_29_LC_22_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_29_LC_22_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_29_LC_22_25_3  (
            .in0(N__39334),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40575),
            .lcout(N_438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_12_LC_22_25_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_12_LC_22_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_12_LC_22_25_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_12_LC_22_25_7  (
            .in0(N__39335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33673),
            .lcout(M_this_oam_ram_write_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_2_LC_22_26_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_2_LC_22_26_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_2_LC_22_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_2_LC_22_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38765),
            .lcout(M_this_scroll_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40455),
            .ce(N__33640),
            .sr(N__39776));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_0_LC_22_27_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_0_LC_22_27_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_0_LC_22_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_0_LC_22_27_2  (
            .in0(_gnd_net_),
            .in1(N__33616),
            .in2(_gnd_net_),
            .in3(N__39370),
            .lcout(M_this_oam_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_1_LC_22_27_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_22_27_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_22_27_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_22_27_4 (
            .in0(N__35470),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40461),
            .ce(N__36029),
            .sr(N__39780));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_1_LC_22_27_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_1_LC_22_27_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_1_LC_22_27_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_1_LC_22_27_5  (
            .in0(N__39371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33598),
            .lcout(M_this_oam_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_25_LC_22_27_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_25_LC_22_27_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_25_LC_22_27_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_25_LC_22_27_6  (
            .in0(N__35471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39369),
            .lcout(N_434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_23_9_6  (
            .in0(N__33571),
            .in1(N__33562),
            .in2(_gnd_net_),
            .in3(N__38900),
            .lcout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_11_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_11_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_spr_ram.mem_mem_7_0_wclke_3_LC_23_11_6  (
            .in0(N__37373),
            .in1(N__37303),
            .in2(N__37474),
            .in3(N__37550),
            .lcout(\this_spr_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_7_LC_23_14_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_7_LC_23_14_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_7_LC_23_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_7_LC_23_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34186),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40366),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_hoffset_q_RNI91DA2_0_LC_23_15_5 .C_ON=1'b0;
    defparam \this_ppu.M_hoffset_q_RNI91DA2_0_LC_23_15_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_hoffset_q_RNI91DA2_0_LC_23_15_5 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_hoffset_q_RNI91DA2_0_LC_23_15_5  (
            .in0(N__34977),
            .in1(N__34158),
            .in2(N__34159),
            .in3(N__35781),
            .lcout(M_this_ppu_spr_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_23_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_23_16_1 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_0_LC_23_16_1  (
            .in0(N__37194),
            .in1(N__35623),
            .in2(N__41056),
            .in3(N__36688),
            .lcout(M_this_spr_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_2_LC_23_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_2_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_2_LC_23_16_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_2_LC_23_16_5  (
            .in0(N__36986),
            .in1(N__37074),
            .in2(_gnd_net_),
            .in3(N__36830),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_3_LC_23_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_3_LC_23_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_3_LC_23_16_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0_3_LC_23_16_7  (
            .in0(N__36987),
            .in1(N__37075),
            .in2(_gnd_net_),
            .in3(N__36831),
            .lcout(\this_ppu.M_this_state_q_srsts_0_i_0_a2_0_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_23_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_23_17_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_ppu.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_23_17_0  (
            .in0(N__36829),
            .in1(N__41259),
            .in2(N__36919),
            .in3(N__33745),
            .lcout(M_this_state_d_0_sqmuxa_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_1_LC_23_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_1_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_i_0_a2_1_1_LC_23_17_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_i_0_a2_1_1_LC_23_17_2  (
            .in0(N__36875),
            .in1(N__33714),
            .in2(N__39920),
            .in3(N__33746),
            .lcout(\this_ppu.N_510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_this_state_q_4_i_0_a2_0_a2_0_LC_23_17_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_4_i_0_a2_0_a2_0_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_4_i_0_a2_0_a2_0_LC_23_17_6 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \this_ppu.un1_M_this_state_q_4_i_0_a2_0_a2_0_LC_23_17_6  (
            .in0(N__33747),
            .in1(N__36967),
            .in2(N__37076),
            .in3(N__33713),
            .lcout(N_608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIPMBQ1_16_LC_23_18_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIPMBQ1_16_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIPMBQ1_16_LC_23_18_0 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIPMBQ1_16_LC_23_18_0  (
            .in0(N__34968),
            .in1(N__35400),
            .in2(_gnd_net_),
            .in3(N__34858),
            .lcout(M_this_ppu_spr_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_15_LC_23_18_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_15_LC_23_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_15_LC_23_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_15_LC_23_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34588),
            .lcout(\this_ppu.un1_M_hoffset_q_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40406),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_14_LC_23_18_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_14_LC_23_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_14_LC_23_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_14_LC_23_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34576),
            .lcout(\this_ppu.un1_M_hoffset_q_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40406),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_23_19_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_23_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_23_19_1  (
            .in0(_gnd_net_),
            .in1(N__41554),
            .in2(_gnd_net_),
            .in3(N__34564),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_23_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_23_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_23_19_3  (
            .in0(_gnd_net_),
            .in1(N__41553),
            .in2(_gnd_net_),
            .in3(N__34501),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_0_14_LC_23_19_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_0_14_LC_23_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI3DGK1_0_14_LC_23_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI3DGK1_0_14_LC_23_19_4  (
            .in0(N__35106),
            .in1(N__35061),
            .in2(N__34423),
            .in3(N__35226),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_c7 ),
            .ltout(\this_ppu.un1_M_oam_cache_read_data_c7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNO_LC_23_19_5 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNO_LC_23_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNO_LC_23_19_5 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNO_LC_23_19_5  (
            .in0(_gnd_net_),
            .in1(N__34342),
            .in2(N__34309),
            .in3(N__34301),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNO_LC_23_19_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNO_LC_23_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNO_LC_23_19_6 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNO_LC_23_19_6  (
            .in0(N__36568),
            .in1(N__35832),
            .in2(N__35338),
            .in3(N__35762),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_2_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_12_LC_23_19_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_12_LC_23_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_12_LC_23_19_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_ppu.oam_cache.read_data_12_LC_23_19_7  (
            .in0(_gnd_net_),
            .in1(N__35350),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.un1_M_hoffset_q_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40416),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNO_LC_23_20_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNO_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNO_LC_23_20_0 .LUT_INIT=16'b0000010111111010;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNO_LC_23_20_0  (
            .in0(N__35750),
            .in1(N__35334),
            .in2(N__35836),
            .in3(N__36562),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_9_LC_23_20_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_9_LC_23_20_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_9_LC_23_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_9_LC_23_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35266),
            .lcout(\this_ppu.un1_M_hoffset_q_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40424),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_8_LC_23_20_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_8_LC_23_20_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_8_LC_23_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_8_LC_23_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35254),
            .lcout(\this_ppu.un1_M_hoffset_q_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40424),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_13_LC_23_20_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_13_LC_23_20_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_13_LC_23_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_13_LC_23_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35242),
            .lcout(\this_ppu.un1_M_hoffset_q_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40424),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI80ET_0_11_LC_23_20_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI80ET_0_11_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI80ET_0_11_LC_23_20_5 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI80ET_0_11_LC_23_20_5  (
            .in0(N__36560),
            .in1(N__35820),
            .in2(N__35923),
            .in3(N__35749),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_c4 ),
            .ltout(\this_ppu.un1_M_oam_cache_read_data_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNO_LC_23_20_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNO_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNO_LC_23_20_6 .LUT_INIT=16'b1100001100110011;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNO_LC_23_20_6  (
            .in0(N__35192),
            .in1(N__35107),
            .in2(N__35080),
            .in3(N__35064),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI80ET_11_LC_23_20_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI80ET_11_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI80ET_11_LC_23_20_7 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI80ET_11_LC_23_20_7  (
            .in0(N__36561),
            .in1(N__35824),
            .in2(N__35924),
            .in3(N__35751),
            .lcout(\this_ppu.read_data_RNI80ET_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_23_21_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_23_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_23_21_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_23_21_0  (
            .in0(N__41468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35002),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_11_LC_23_21_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_11_LC_23_21_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_11_LC_23_21_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_11_LC_23_21_1  (
            .in0(N__35941),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.un1_M_hoffset_q_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40432),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNO_LC_23_21_3 .C_ON=1'b0;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNO_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNO_LC_23_21_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNO_LC_23_21_3  (
            .in0(N__35899),
            .in1(N__35825),
            .in2(_gnd_net_),
            .in3(N__35752),
            .lcout(\this_ppu.un1_M_oam_cache_read_data_3_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_4_c5_LC_23_21_5 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_4_c5_LC_23_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_4_c5_LC_23_21_5 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \this_ppu.un1_oam_data_1_4_c5_LC_23_21_5  (
            .in0(N__38566),
            .in1(N__38443),
            .in2(N__38512),
            .in3(N__38359),
            .lcout(\this_ppu.un1_oam_data_1_4_c5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_23_21_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_23_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_23_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_23_21_7  (
            .in0(_gnd_net_),
            .in1(N__41469),
            .in2(_gnd_net_),
            .in3(N__35679),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_14_LC_23_22_0.C_ON=1'b0;
    defparam M_this_ext_address_q_14_LC_23_22_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_14_LC_23_22_0.LUT_INIT=16'b1101100011001100;
    LogicCell40 M_this_ext_address_q_14_LC_23_22_0 (
            .in0(N__40717),
            .in1(N__37984),
            .in2(N__36308),
            .in3(N__40887),
            .lcout(M_this_ext_address_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40441),
            .ce(),
            .sr(N__39762));
    defparam M_this_ext_address_q_8_LC_23_22_1.C_ON=1'b0;
    defparam M_this_ext_address_q_8_LC_23_22_1.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_8_LC_23_22_1.LUT_INIT=16'b1111110100100000;
    LogicCell40 M_this_ext_address_q_8_LC_23_22_1 (
            .in0(N__40885),
            .in1(N__40719),
            .in2(N__35618),
            .in3(N__37810),
            .lcout(M_this_ext_address_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40441),
            .ce(),
            .sr(N__39762));
    defparam M_this_ext_address_q_9_LC_23_22_2.C_ON=1'b0;
    defparam M_this_ext_address_q_9_LC_23_22_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_9_LC_23_22_2.LUT_INIT=16'b1111010010110000;
    LogicCell40 M_this_ext_address_q_9_LC_23_22_2 (
            .in0(N__40718),
            .in1(N__40886),
            .in2(N__37777),
            .in3(N__35498),
            .lcout(M_this_ext_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40441),
            .ce(),
            .sr(N__39762));
    defparam \this_ppu.oam_cache.read_data_16_LC_23_23_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_16_LC_23_23_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_16_LC_23_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_16_LC_23_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35413),
            .lcout(\this_ppu.M_oam_cache_read_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40446),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_20_LC_23_23_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_20_LC_23_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_20_LC_23_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_20_LC_23_23_6  (
            .in0(_gnd_net_),
            .in1(N__35380),
            .in2(_gnd_net_),
            .in3(N__39314),
            .lcout(M_this_oam_ram_write_data_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_6_LC_23_24_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_23_24_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_23_24_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_23_24_1 (
            .in0(N__36309),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40451),
            .ce(N__36030),
            .sr(N__39766));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_7_LC_23_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_7_LC_23_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_7_LC_23_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_7_LC_23_24_2  (
            .in0(_gnd_net_),
            .in1(N__36073),
            .in2(_gnd_net_),
            .in3(N__39315),
            .lcout(M_this_oam_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_7_LC_23_24_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_23_24_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_23_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_23_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36477),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40451),
            .ce(N__36030),
            .sr(N__39766));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_3_LC_23_25_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_3_LC_23_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_3_LC_23_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_3_LC_23_25_0  (
            .in0(_gnd_net_),
            .in1(N__36055),
            .in2(_gnd_net_),
            .in3(N__39316),
            .lcout(M_this_oam_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_3_LC_23_25_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_23_25_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_23_25_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_23_25_1 (
            .in0(N__39478),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40456),
            .ce(N__36031),
            .sr(N__39771));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_4_LC_23_25_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_4_LC_23_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_4_LC_23_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_4_LC_23_25_3  (
            .in0(N__39317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36037),
            .lcout(M_this_oam_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_4_LC_23_25_4.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_23_25_4.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_23_25_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_23_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41029),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40456),
            .ce(N__36031),
            .sr(N__39771));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_23_LC_23_26_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_23_LC_23_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_23_LC_23_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_23_LC_23_26_3  (
            .in0(_gnd_net_),
            .in1(N__35974),
            .in2(_gnd_net_),
            .in3(N__39318),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_23_26_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_23_26_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_23_26_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_23_26_6  (
            .in0(_gnd_net_),
            .in1(N__41584),
            .in2(_gnd_net_),
            .in3(N__39102),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_31_LC_23_27_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_31_LC_23_27_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_31_LC_23_27_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_31_LC_23_27_1  (
            .in0(_gnd_net_),
            .in1(N__36486),
            .in2(_gnd_net_),
            .in3(N__39308),
            .lcout(N_440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_28_LC_23_27_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_28_LC_23_27_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_28_LC_23_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_28_LC_23_27_4  (
            .in0(_gnd_net_),
            .in1(N__40983),
            .in2(_gnd_net_),
            .in3(N__39307),
            .lcout(N_437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_22_LC_23_28_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_22_LC_23_28_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_22_LC_23_28_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_22_LC_23_28_3  (
            .in0(_gnd_net_),
            .in1(N__36331),
            .in2(_gnd_net_),
            .in3(N__39313),
            .lcout(M_this_oam_ram_write_data_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_30_LC_23_28_5 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_30_LC_23_28_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_30_LC_23_28_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_30_LC_23_28_5  (
            .in0(_gnd_net_),
            .in1(N__36313),
            .in2(_gnd_net_),
            .in3(N__39312),
            .lcout(N_439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_9_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_9_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_9_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_spr_ram.mem_mem_6_0_wclke_3_LC_24_9_3  (
            .in0(N__37384),
            .in1(N__37476),
            .in2(N__37305),
            .in3(N__37555),
            .lcout(\this_spr_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_11_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_11_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_spr_ram.mem_mem_5_0_wclke_3_LC_24_11_3  (
            .in0(N__37379),
            .in1(N__37467),
            .in2(N__37306),
            .in3(N__37551),
            .lcout(\this_spr_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_24_11_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_24_11_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_24_11_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_24_11_5  (
            .in0(N__36145),
            .in1(N__36139),
            .in2(_gnd_net_),
            .in3(N__38899),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_13_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_13_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_spr_ram.mem_mem_0_0_wclke_3_LC_24_13_0  (
            .in0(N__37301),
            .in1(N__37375),
            .in2(N__37475),
            .in3(N__37547),
            .lcout(\this_spr_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_13_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_spr_ram.mem_mem_1_0_wclke_3_LC_24_13_3  (
            .in0(N__37548),
            .in1(N__37466),
            .in2(N__37383),
            .in3(N__37302),
            .lcout(\this_spr_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_24_14_3 .C_ON=1'b0;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_24_14_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_24_14_3 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \this_ppu.M_this_spr_ram_write_data_1_0_i_3_LC_24_14_3  (
            .in0(N__36429),
            .in1(N__37201),
            .in2(N__39516),
            .in3(N__36679),
            .lcout(M_this_spr_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_1_3_LC_24_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_1_3_LC_24_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_i_0_a2_1_3_LC_24_16_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_i_0_a2_1_3_LC_24_16_0  (
            .in0(N__37063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36988),
            .lcout(\this_ppu.N_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_24_17_5.C_ON=1'b0;
    defparam M_this_substate_q_LC_24_17_5.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_24_17_5.LUT_INIT=16'b1010110011001100;
    LogicCell40 M_this_substate_q_LC_24_17_5 (
            .in0(N__36910),
            .in1(N__36832),
            .in2(N__36894),
            .in3(N__36844),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40407),
            .ce(),
            .sr(N__39754));
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_i_LC_24_19_0 .C_ON=1'b0;
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_i_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_this_state_q_1_i_0_0_i_LC_24_19_0 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \this_ppu.un1_M_this_state_q_1_i_0_0_i_LC_24_19_0  (
            .in0(N__36810),
            .in1(N__36738),
            .in2(N__36687),
            .in3(N__40855),
            .lcout(N_312_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_10_LC_24_19_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_10_LC_24_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_10_LC_24_19_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \this_ppu.oam_cache.read_data_10_LC_24_19_4  (
            .in0(_gnd_net_),
            .in1(N__36595),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.un1_M_hoffset_q_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40425),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_24_19_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_24_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_24_19_7  (
            .in0(_gnd_net_),
            .in1(N__41602),
            .in2(_gnd_net_),
            .in3(N__38442),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_15_LC_24_20_0.C_ON=1'b0;
    defparam M_this_ext_address_q_15_LC_24_20_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_15_LC_24_20_0.LUT_INIT=16'b1111110100001000;
    LogicCell40 M_this_ext_address_q_15_LC_24_20_0 (
            .in0(N__40879),
            .in1(N__36476),
            .in2(N__40720),
            .in3(N__37945),
            .lcout(M_this_ext_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam M_this_ctrl_flags_q_7_LC_24_20_1.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_7_LC_24_20_1.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_7_LC_24_20_1.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_this_ctrl_flags_q_7_LC_24_20_1 (
            .in0(N__37743),
            .in1(N__36523),
            .in2(N__36485),
            .in3(N__40882),
            .lcout(M_this_ctrl_flags_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam M_this_ext_address_q_0_LC_24_20_4.C_ON=1'b0;
    defparam M_this_ext_address_q_0_LC_24_20_4.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_0_LC_24_20_4.LUT_INIT=16'b0011000111000100;
    LogicCell40 M_this_ext_address_q_0_LC_24_20_4 (
            .in0(N__40880),
            .in1(N__37700),
            .in2(N__40721),
            .in3(N__37731),
            .lcout(M_this_ext_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam M_this_ext_address_q_1_LC_24_20_5.C_ON=1'b0;
    defparam M_this_ext_address_q_1_LC_24_20_5.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_1_LC_24_20_5.LUT_INIT=16'b0101101000010010;
    LogicCell40 M_this_ext_address_q_1_LC_24_20_5 (
            .in0(N__37668),
            .in1(N__40883),
            .in2(N__37651),
            .in3(N__40699),
            .lcout(M_this_ext_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam M_this_ext_address_q_2_LC_24_20_6.C_ON=1'b0;
    defparam M_this_ext_address_q_2_LC_24_20_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_2_LC_24_20_6.LUT_INIT=16'b0011000111000100;
    LogicCell40 M_this_ext_address_q_2_LC_24_20_6 (
            .in0(N__40881),
            .in1(N__37626),
            .in2(N__40722),
            .in3(N__37609),
            .lcout(M_this_ext_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam M_this_ext_address_q_3_LC_24_20_7.C_ON=1'b0;
    defparam M_this_ext_address_q_3_LC_24_20_7.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_3_LC_24_20_7.LUT_INIT=16'b0101101000010010;
    LogicCell40 M_this_ext_address_q_3_LC_24_20_7 (
            .in0(N__37584),
            .in1(N__40884),
            .in2(N__37567),
            .in3(N__40700),
            .lcout(M_this_ext_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40433),
            .ce(),
            .sr(N__39755));
    defparam un1_M_this_ext_address_q_cry_0_c_LC_24_21_0.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_0_c_LC_24_21_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_0_c_LC_24_21_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_ext_address_q_cry_0_c_LC_24_21_0 (
            .in0(_gnd_net_),
            .in1(N__37732),
            .in2(N__37704),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_24_21_0_),
            .carryout(un1_M_this_ext_address_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_24_21_1.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_24_21_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_24_21_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_0_THRU_LUT4_0_LC_24_21_1 (
            .in0(_gnd_net_),
            .in1(N__37667),
            .in2(_gnd_net_),
            .in3(N__37639),
            .lcout(un1_M_this_ext_address_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_0),
            .carryout(un1_M_this_ext_address_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_24_21_2.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_24_21_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_24_21_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_1_THRU_LUT4_0_LC_24_21_2 (
            .in0(_gnd_net_),
            .in1(N__37625),
            .in2(_gnd_net_),
            .in3(N__37603),
            .lcout(un1_M_this_ext_address_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_1),
            .carryout(un1_M_this_ext_address_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_24_21_3.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_24_21_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_24_21_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_2_THRU_LUT4_0_LC_24_21_3 (
            .in0(_gnd_net_),
            .in1(N__37583),
            .in2(_gnd_net_),
            .in3(N__37558),
            .lcout(un1_M_this_ext_address_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_2),
            .carryout(un1_M_this_ext_address_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_24_21_4.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_24_21_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_24_21_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_3_THRU_LUT4_0_LC_24_21_4 (
            .in0(_gnd_net_),
            .in1(N__38625),
            .in2(_gnd_net_),
            .in3(N__37849),
            .lcout(un1_M_this_ext_address_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_3),
            .carryout(un1_M_this_ext_address_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_24_21_5.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_24_21_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_24_21_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_4_THRU_LUT4_0_LC_24_21_5 (
            .in0(_gnd_net_),
            .in1(N__41229),
            .in2(_gnd_net_),
            .in3(N__37846),
            .lcout(un1_M_this_ext_address_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_4),
            .carryout(un1_M_this_ext_address_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_24_21_6.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_24_21_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_24_21_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_5_THRU_LUT4_0_LC_24_21_6 (
            .in0(_gnd_net_),
            .in1(N__41184),
            .in2(_gnd_net_),
            .in3(N__37843),
            .lcout(un1_M_this_ext_address_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_5),
            .carryout(un1_M_this_ext_address_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_24_21_7.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_24_21_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_24_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_M_this_ext_address_q_cry_6_THRU_LUT4_0_LC_24_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41136),
            .in3(N__37840),
            .lcout(un1_M_this_ext_address_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_6),
            .carryout(un1_M_this_ext_address_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_24_22_0.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_24_22_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_24_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_7_c_RNIQ14F_LC_24_22_0 (
            .in0(_gnd_net_),
            .in1(N__37821),
            .in2(_gnd_net_),
            .in3(N__37804),
            .lcout(un1_M_this_ext_address_q_cry_7_c_RNIQ14FZ0),
            .ltout(),
            .carryin(bfn_24_22_0_),
            .carryout(un1_M_this_ext_address_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_24_22_1.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_24_22_1.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_24_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_8_c_RNIS45F_LC_24_22_1 (
            .in0(_gnd_net_),
            .in1(N__37788),
            .in2(_gnd_net_),
            .in3(N__37765),
            .lcout(un1_M_this_ext_address_q_cry_8_c_RNIS45FZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_8),
            .carryout(un1_M_this_ext_address_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_24_22_2.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_24_22_2.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_24_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_9_c_RNI55NH_LC_24_22_2 (
            .in0(_gnd_net_),
            .in1(N__38652),
            .in2(_gnd_net_),
            .in3(N__37762),
            .lcout(un1_M_this_ext_address_q_cry_9_c_RNI55NHZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_9),
            .carryout(un1_M_this_ext_address_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_24_22_3.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_24_22_3.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_24_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_10_c_RNIEGOA_LC_24_22_3 (
            .in0(_gnd_net_),
            .in1(N__41082),
            .in2(_gnd_net_),
            .in3(N__37759),
            .lcout(un1_M_this_ext_address_q_cry_10_c_RNIEGOAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_10),
            .carryout(un1_M_this_ext_address_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_24_22_4.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_24_22_4.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_24_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_M_this_ext_address_q_cry_11_c_RNIGJPA_LC_24_22_4 (
            .in0(_gnd_net_),
            .in1(N__40929),
            .in2(_gnd_net_),
            .in3(N__37756),
            .lcout(un1_M_this_ext_address_q_cry_11_c_RNIGJPAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_11),
            .carryout(un1_M_this_ext_address_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_24_22_5.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_24_22_5.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_24_22_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_ext_address_q_cry_12_c_RNIIMQA_LC_24_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40488),
            .in3(N__38014),
            .lcout(un1_M_this_ext_address_q_cry_12_c_RNIIMQAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_12),
            .carryout(un1_M_this_ext_address_q_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_24_22_6.C_ON=1'b1;
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_24_22_6.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_24_22_6.LUT_INIT=16'b1010010101011010;
    LogicCell40 un1_M_this_ext_address_q_cry_13_c_RNIKPRA_LC_24_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38001),
            .in3(N__37978),
            .lcout(un1_M_this_ext_address_q_cry_13_c_RNIKPRAZ0),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_13),
            .carryout(un1_M_this_ext_address_q_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_24_22_7.C_ON=1'b0;
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_24_22_7.SEQ_MODE=4'b0000;
    defparam un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_24_22_7.LUT_INIT=16'b0101010110101010;
    LogicCell40 un1_M_this_ext_address_q_cry_14_c_RNIMSSA_LC_24_22_7 (
            .in0(N__37965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37948),
            .lcout(un1_M_this_ext_address_q_cry_14_c_RNIMSSAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_24_23_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_24_23_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_24_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_24_23_1  (
            .in0(_gnd_net_),
            .in1(N__37936),
            .in2(_gnd_net_),
            .in3(N__41564),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_24_23_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_24_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_24_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_24_23_3  (
            .in0(_gnd_net_),
            .in1(N__37918),
            .in2(_gnd_net_),
            .in3(N__41565),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_24_23_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_24_23_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_24_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_24_23_4  (
            .in0(N__38236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41568),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_24_23_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_24_23_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_24_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_24_23_5  (
            .in0(_gnd_net_),
            .in1(N__37891),
            .in2(_gnd_net_),
            .in3(N__41566),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_24_23_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_24_23_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_24_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_24_23_6  (
            .in0(_gnd_net_),
            .in1(N__41569),
            .in2(_gnd_net_),
            .in3(N__39056),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_24_23_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_24_23_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_24_23_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_24_23_7  (
            .in0(_gnd_net_),
            .in1(N__37867),
            .in2(_gnd_net_),
            .in3(N__41567),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_24_24_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_24_24_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_24_24_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_24_24_0  (
            .in0(N__41574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38149),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_24_24_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_24_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_24_24_1  (
            .in0(_gnd_net_),
            .in1(N__41575),
            .in2(_gnd_net_),
            .in3(N__38131),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_10_LC_24_24_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_10_LC_24_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_10_LC_24_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_10_LC_24_24_2  (
            .in0(_gnd_net_),
            .in1(N__38113),
            .in2(_gnd_net_),
            .in3(N__39375),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_6_LC_24_24_4 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_6_LC_24_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_6_LC_24_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_6_LC_24_24_4  (
            .in0(_gnd_net_),
            .in1(N__38095),
            .in2(_gnd_net_),
            .in3(N__39377),
            .lcout(M_this_oam_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_11_LC_24_24_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_11_LC_24_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_11_LC_24_24_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_11_LC_24_24_6  (
            .in0(_gnd_net_),
            .in1(N__38080),
            .in2(_gnd_net_),
            .in3(N__39376),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_24_24_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_24_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_24_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_24_24_7  (
            .in0(_gnd_net_),
            .in1(N__41573),
            .in2(_gnd_net_),
            .in3(N__38260),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un12lto7_4_LC_24_25_0 .C_ON=1'b0;
    defparam \this_ppu.un12lto7_4_LC_24_25_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un12lto7_4_LC_24_25_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un12lto7_4_LC_24_25_0  (
            .in0(N__38319),
            .in1(N__38340),
            .in2(N__38302),
            .in3(N__38034),
            .lcout(\this_ppu.un12lto7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_24_25_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_24_25_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_24_25_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_24_25_1  (
            .in0(N__38035),
            .in1(_gnd_net_),
            .in2(N__41603),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_24_25_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_24_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_24_25_2  (
            .in0(_gnd_net_),
            .in1(N__41580),
            .in2(_gnd_net_),
            .in3(N__38341),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_24_25_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_24_25_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_24_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_24_25_3  (
            .in0(N__41581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38320),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_24_25_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_24_25_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_24_25_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_24_25_4  (
            .in0(N__38301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41582),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_24_25_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_24_25_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_24_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_24_25_5  (
            .in0(N__41583),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38218),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_24_25_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_24_25_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_24_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_24_25_6  (
            .in0(N__38245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41576),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un12lto7_5_LC_24_25_7 .C_ON=1'b0;
    defparam \this_ppu.un12lto7_5_LC_24_25_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un12lto7_5_LC_24_25_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un12lto7_5_LC_24_25_7  (
            .in0(N__38256),
            .in1(N__38244),
            .in2(N__38235),
            .in3(N__38217),
            .lcout(\this_ppu.un12lto7Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_24_26_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_24_26_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_24_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_24_26_0  (
            .in0(_gnd_net_),
            .in1(N__38200),
            .in2(_gnd_net_),
            .in3(N__41585),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNO_LC_24_26_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNO_LC_24_26_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNO_LC_24_26_1 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_3_c_RNO_LC_24_26_1  (
            .in0(N__38430),
            .in1(N__39092),
            .in2(N__38563),
            .in3(N__39046),
            .lcout(\this_ppu.un1_oam_data_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_24_26_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_24_26_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_24_26_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_24_26_2  (
            .in0(_gnd_net_),
            .in1(N__38167),
            .in2(_gnd_net_),
            .in3(N__41586),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNO_LC_24_26_3 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNO_LC_24_26_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNO_LC_24_26_3 .LUT_INIT=16'b1001001111000011;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_4_c_RNO_LC_24_26_3  (
            .in0(N__38431),
            .in1(N__38500),
            .in2(N__38564),
            .in3(N__38355),
            .lcout(\this_ppu.un1_oam_data_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_24_26_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_24_26_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_24_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_24_26_4  (
            .in0(_gnd_net_),
            .in1(N__38581),
            .in2(_gnd_net_),
            .in3(N__41587),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_24_26_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_24_26_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_24_26_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_24_26_5  (
            .in0(N__38556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41589),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_24_26_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_24_26_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_24_26_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_24_26_6  (
            .in0(N__38501),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41588),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_24_26_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_24_26_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_24_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_24_26_7  (
            .in0(_gnd_net_),
            .in1(N__38461),
            .in2(_gnd_net_),
            .in3(N__41590),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNO_LC_24_27_1 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNO_LC_24_27_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_RNO_LC_24_27_1 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_2_c_RNO_LC_24_27_1  (
            .in0(N__38415),
            .in1(N__39083),
            .in2(_gnd_net_),
            .in3(N__39034),
            .lcout(\this_ppu.un1_oam_data_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_17_LC_24_27_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_17_LC_24_27_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_0_a2_17_LC_24_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_0_a2_17_LC_24_27_2  (
            .in0(_gnd_net_),
            .in1(N__38374),
            .in2(_gnd_net_),
            .in3(N__39374),
            .lcout(M_this_oam_ram_write_data_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_4_ac0_1_LC_24_27_3 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_4_ac0_1_LC_24_27_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_4_ac0_1_LC_24_27_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.un1_oam_data_1_4_ac0_1_LC_24_27_3  (
            .in0(_gnd_net_),
            .in1(N__39081),
            .in2(_gnd_net_),
            .in3(N__39032),
            .lcout(\this_ppu.un1_oam_data_1_4_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_24_27_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_24_27_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_24_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_24_27_4  (
            .in0(N__41592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39154),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_24_27_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_24_27_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_24_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_24_27_5  (
            .in0(_gnd_net_),
            .in1(N__41591),
            .in2(_gnd_net_),
            .in3(N__39133),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_26_LC_24_27_6 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_26_LC_24_27_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_26_LC_24_27_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_26_LC_24_27_6  (
            .in0(N__38754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39373),
            .lcout(N_435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_1_c_RNO_LC_24_27_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_RNO_LC_24_27_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_RNO_LC_24_27_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_1_c_RNO_LC_24_27_7  (
            .in0(_gnd_net_),
            .in1(N__39082),
            .in2(_gnd_net_),
            .in3(N__39033),
            .lcout(\this_ppu.un1_oam_data_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_26_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_26_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_26_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_26_9_6  (
            .in0(N__38998),
            .in1(N__38992),
            .in2(_gnd_net_),
            .in3(N__38929),
            .lcout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_26_10_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_26_10_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_26_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_26_10_4  (
            .in0(N__38965),
            .in1(N__38956),
            .in2(_gnd_net_),
            .in3(N__38928),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_10_LC_26_22_0.C_ON=1'b0;
    defparam M_this_ext_address_q_10_LC_26_22_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_10_LC_26_22_0.LUT_INIT=16'b1011100010101010;
    LogicCell40 M_this_ext_address_q_10_LC_26_22_0 (
            .in0(N__38800),
            .in1(N__40710),
            .in2(N__38760),
            .in3(N__40909),
            .lcout(M_this_ext_address_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_4_LC_26_22_1.C_ON=1'b0;
    defparam M_this_ext_address_q_4_LC_26_22_1.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_4_LC_26_22_1.LUT_INIT=16'b0011000111000100;
    LogicCell40 M_this_ext_address_q_4_LC_26_22_1 (
            .in0(N__40907),
            .in1(N__38615),
            .in2(N__40725),
            .in3(N__38638),
            .lcout(M_this_ext_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_5_LC_26_22_2.C_ON=1'b0;
    defparam M_this_ext_address_q_5_LC_26_22_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_5_LC_26_22_2.LUT_INIT=16'b0110000001100110;
    LogicCell40 M_this_ext_address_q_5_LC_26_22_2 (
            .in0(N__41222),
            .in1(N__41245),
            .in2(N__40723),
            .in3(N__40911),
            .lcout(M_this_ext_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_6_LC_26_22_3.C_ON=1'b0;
    defparam M_this_ext_address_q_6_LC_26_22_3.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_6_LC_26_22_3.LUT_INIT=16'b0011000111000100;
    LogicCell40 M_this_ext_address_q_6_LC_26_22_3 (
            .in0(N__40908),
            .in1(N__41177),
            .in2(N__40726),
            .in3(N__41203),
            .lcout(M_this_ext_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_7_LC_26_22_4.C_ON=1'b0;
    defparam M_this_ext_address_q_7_LC_26_22_4.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_7_LC_26_22_4.LUT_INIT=16'b0110000001100110;
    LogicCell40 M_this_ext_address_q_7_LC_26_22_4 (
            .in0(N__41120),
            .in1(N__41158),
            .in2(N__40724),
            .in3(N__40912),
            .lcout(M_this_ext_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_11_LC_26_22_5.C_ON=1'b0;
    defparam M_this_ext_address_q_11_LC_26_22_5.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_11_LC_26_22_5.LUT_INIT=16'b1111110100100000;
    LogicCell40 M_this_ext_address_q_11_LC_26_22_5 (
            .in0(N__40905),
            .in1(N__40702),
            .in2(N__39505),
            .in3(N__41101),
            .lcout(M_this_ext_address_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_12_LC_26_22_6.C_ON=1'b0;
    defparam M_this_ext_address_q_12_LC_26_22_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_12_LC_26_22_6.LUT_INIT=16'b1101100011001100;
    LogicCell40 M_this_ext_address_q_12_LC_26_22_6 (
            .in0(N__40701),
            .in1(N__41065),
            .in2(N__41040),
            .in3(N__40910),
            .lcout(M_this_ext_address_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam M_this_ext_address_q_13_LC_26_22_7.C_ON=1'b0;
    defparam M_this_ext_address_q_13_LC_26_22_7.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_13_LC_26_22_7.LUT_INIT=16'b1111110100100000;
    LogicCell40 M_this_ext_address_q_13_LC_26_22_7 (
            .in0(N__40906),
            .in1(N__40703),
            .in2(N__40582),
            .in3(N__40501),
            .lcout(M_this_ext_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40459),
            .ce(),
            .sr(N__39756));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_26_23_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_26_23_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_26_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_26_23_3  (
            .in0(_gnd_net_),
            .in1(N__39538),
            .in2(_gnd_net_),
            .in3(N__41597),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_27_LC_26_29_2 .C_ON=1'b0;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_27_LC_26_29_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_oam_ram_write_data_i_i_a2_27_LC_26_29_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.M_this_oam_ram_write_data_i_i_a2_27_LC_26_29_2  (
            .in0(N__39440),
            .in1(N__39319),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_27_27_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_27_27_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_27_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_27_27_2  (
            .in0(_gnd_net_),
            .in1(N__41638),
            .in2(_gnd_net_),
            .in3(N__41605),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_28_24_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_28_24_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_28_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_28_24_2  (
            .in0(_gnd_net_),
            .in1(N__41617),
            .in2(_gnd_net_),
            .in3(N__41604),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1_0_LC_31_28_1 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1_0_LC_31_28_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1_0_LC_31_28_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1_0_LC_31_28_1  (
            .in0(N__41344),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41326),
            .lcout(\this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_0_LC_32_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_0_LC_32_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_0_LC_32_17_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_this_state_q_srsts_0_o2_0_i_a2_0_0_LC_32_17_7  (
            .in0(N__41317),
            .in1(N__41311),
            .in2(N__41299),
            .in3(N__41284),
            .lcout(\this_ppu.N_173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cu_top_0
