// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec 10 2020 17:46:48

// File Generated:     Jun 1 2022 00:08:23

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cu_top_0" view "INTERFACE"

module cu_top_0 (
    port_address,
    port_data,
    debug,
    rgb,
    led,
    vsync,
    vblank,
    rst_n,
    port_rw,
    port_nmib,
    port_enb,
    port_dmab,
    port_data_rw,
    port_clk,
    hsync,
    hblank,
    clk);

    inout [15:0] port_address;
    input [7:0] port_data;
    output [1:0] debug;
    output [5:0] rgb;
    output [7:0] led;
    output vsync;
    output vblank;
    input rst_n;
    inout port_rw;
    output port_nmib;
    input port_enb;
    output port_dmab;
    output port_data_rw;
    input port_clk;
    output hsync;
    output hblank;
    input clk;

    wire N__40097;
    wire N__40096;
    wire N__40095;
    wire N__40086;
    wire N__40085;
    wire N__40084;
    wire N__40077;
    wire N__40076;
    wire N__40075;
    wire N__40068;
    wire N__40067;
    wire N__40066;
    wire N__40059;
    wire N__40058;
    wire N__40057;
    wire N__40050;
    wire N__40049;
    wire N__40048;
    wire N__40041;
    wire N__40040;
    wire N__40039;
    wire N__40032;
    wire N__40031;
    wire N__40030;
    wire N__40023;
    wire N__40022;
    wire N__40021;
    wire N__40014;
    wire N__40013;
    wire N__40012;
    wire N__40005;
    wire N__40004;
    wire N__40003;
    wire N__39996;
    wire N__39995;
    wire N__39994;
    wire N__39987;
    wire N__39986;
    wire N__39985;
    wire N__39978;
    wire N__39977;
    wire N__39976;
    wire N__39969;
    wire N__39968;
    wire N__39967;
    wire N__39960;
    wire N__39959;
    wire N__39958;
    wire N__39951;
    wire N__39950;
    wire N__39949;
    wire N__39942;
    wire N__39941;
    wire N__39940;
    wire N__39933;
    wire N__39932;
    wire N__39931;
    wire N__39924;
    wire N__39923;
    wire N__39922;
    wire N__39915;
    wire N__39914;
    wire N__39913;
    wire N__39906;
    wire N__39905;
    wire N__39904;
    wire N__39897;
    wire N__39896;
    wire N__39895;
    wire N__39888;
    wire N__39887;
    wire N__39886;
    wire N__39879;
    wire N__39878;
    wire N__39877;
    wire N__39870;
    wire N__39869;
    wire N__39868;
    wire N__39861;
    wire N__39860;
    wire N__39859;
    wire N__39852;
    wire N__39851;
    wire N__39850;
    wire N__39843;
    wire N__39842;
    wire N__39841;
    wire N__39834;
    wire N__39833;
    wire N__39832;
    wire N__39825;
    wire N__39824;
    wire N__39823;
    wire N__39816;
    wire N__39815;
    wire N__39814;
    wire N__39807;
    wire N__39806;
    wire N__39805;
    wire N__39798;
    wire N__39797;
    wire N__39796;
    wire N__39789;
    wire N__39788;
    wire N__39787;
    wire N__39780;
    wire N__39779;
    wire N__39778;
    wire N__39771;
    wire N__39770;
    wire N__39769;
    wire N__39762;
    wire N__39761;
    wire N__39760;
    wire N__39753;
    wire N__39752;
    wire N__39751;
    wire N__39744;
    wire N__39743;
    wire N__39742;
    wire N__39735;
    wire N__39734;
    wire N__39733;
    wire N__39726;
    wire N__39725;
    wire N__39724;
    wire N__39717;
    wire N__39716;
    wire N__39715;
    wire N__39708;
    wire N__39707;
    wire N__39706;
    wire N__39699;
    wire N__39698;
    wire N__39697;
    wire N__39690;
    wire N__39689;
    wire N__39688;
    wire N__39681;
    wire N__39680;
    wire N__39679;
    wire N__39672;
    wire N__39671;
    wire N__39670;
    wire N__39663;
    wire N__39662;
    wire N__39661;
    wire N__39654;
    wire N__39653;
    wire N__39652;
    wire N__39645;
    wire N__39644;
    wire N__39643;
    wire N__39636;
    wire N__39635;
    wire N__39634;
    wire N__39617;
    wire N__39614;
    wire N__39611;
    wire N__39608;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39593;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39581;
    wire N__39578;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39538;
    wire N__39533;
    wire N__39530;
    wire N__39527;
    wire N__39526;
    wire N__39525;
    wire N__39524;
    wire N__39523;
    wire N__39522;
    wire N__39521;
    wire N__39520;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39514;
    wire N__39509;
    wire N__39500;
    wire N__39491;
    wire N__39488;
    wire N__39481;
    wire N__39478;
    wire N__39475;
    wire N__39472;
    wire N__39469;
    wire N__39464;
    wire N__39461;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39434;
    wire N__39433;
    wire N__39432;
    wire N__39431;
    wire N__39430;
    wire N__39429;
    wire N__39428;
    wire N__39427;
    wire N__39426;
    wire N__39425;
    wire N__39424;
    wire N__39423;
    wire N__39422;
    wire N__39421;
    wire N__39420;
    wire N__39419;
    wire N__39418;
    wire N__39417;
    wire N__39416;
    wire N__39415;
    wire N__39414;
    wire N__39413;
    wire N__39412;
    wire N__39411;
    wire N__39410;
    wire N__39409;
    wire N__39408;
    wire N__39407;
    wire N__39406;
    wire N__39405;
    wire N__39404;
    wire N__39403;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39399;
    wire N__39398;
    wire N__39397;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39393;
    wire N__39392;
    wire N__39391;
    wire N__39390;
    wire N__39389;
    wire N__39388;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39384;
    wire N__39383;
    wire N__39382;
    wire N__39381;
    wire N__39380;
    wire N__39379;
    wire N__39378;
    wire N__39377;
    wire N__39376;
    wire N__39375;
    wire N__39374;
    wire N__39373;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39369;
    wire N__39368;
    wire N__39367;
    wire N__39366;
    wire N__39365;
    wire N__39364;
    wire N__39363;
    wire N__39362;
    wire N__39361;
    wire N__39360;
    wire N__39359;
    wire N__39358;
    wire N__39357;
    wire N__39356;
    wire N__39355;
    wire N__39354;
    wire N__39353;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39349;
    wire N__39348;
    wire N__39347;
    wire N__39346;
    wire N__39345;
    wire N__39344;
    wire N__39343;
    wire N__39342;
    wire N__39341;
    wire N__39340;
    wire N__39339;
    wire N__39338;
    wire N__39337;
    wire N__39336;
    wire N__39335;
    wire N__39334;
    wire N__39333;
    wire N__39332;
    wire N__39331;
    wire N__39330;
    wire N__39329;
    wire N__39328;
    wire N__39327;
    wire N__39326;
    wire N__39325;
    wire N__39324;
    wire N__39323;
    wire N__39322;
    wire N__39321;
    wire N__39320;
    wire N__39319;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39313;
    wire N__39312;
    wire N__39311;
    wire N__39310;
    wire N__39309;
    wire N__39308;
    wire N__39307;
    wire N__39306;
    wire N__39305;
    wire N__39304;
    wire N__39303;
    wire N__39302;
    wire N__39301;
    wire N__39300;
    wire N__39299;
    wire N__39298;
    wire N__39297;
    wire N__39296;
    wire N__39295;
    wire N__39294;
    wire N__39293;
    wire N__39292;
    wire N__39291;
    wire N__39290;
    wire N__39289;
    wire N__39288;
    wire N__39287;
    wire N__39286;
    wire N__39285;
    wire N__39284;
    wire N__39283;
    wire N__39282;
    wire N__39281;
    wire N__39280;
    wire N__38969;
    wire N__38966;
    wire N__38963;
    wire N__38962;
    wire N__38961;
    wire N__38960;
    wire N__38959;
    wire N__38958;
    wire N__38957;
    wire N__38956;
    wire N__38955;
    wire N__38954;
    wire N__38953;
    wire N__38952;
    wire N__38951;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38917;
    wire N__38914;
    wire N__38911;
    wire N__38910;
    wire N__38909;
    wire N__38904;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38896;
    wire N__38895;
    wire N__38894;
    wire N__38891;
    wire N__38890;
    wire N__38887;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38874;
    wire N__38871;
    wire N__38868;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38845;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38828;
    wire N__38825;
    wire N__38822;
    wire N__38817;
    wire N__38812;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38780;
    wire N__38777;
    wire N__38774;
    wire N__38773;
    wire N__38770;
    wire N__38769;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38761;
    wire N__38760;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38689;
    wire N__38686;
    wire N__38681;
    wire N__38676;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38641;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38629;
    wire N__38628;
    wire N__38627;
    wire N__38626;
    wire N__38625;
    wire N__38624;
    wire N__38621;
    wire N__38620;
    wire N__38619;
    wire N__38618;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38591;
    wire N__38588;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38578;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38564;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38540;
    wire N__38537;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38519;
    wire N__38516;
    wire N__38513;
    wire N__38510;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38495;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38483;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38465;
    wire N__38462;
    wire N__38459;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38449;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38435;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38396;
    wire N__38393;
    wire N__38392;
    wire N__38389;
    wire N__38386;
    wire N__38383;
    wire N__38378;
    wire N__38375;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38365;
    wire N__38362;
    wire N__38359;
    wire N__38356;
    wire N__38351;
    wire N__38348;
    wire N__38347;
    wire N__38346;
    wire N__38345;
    wire N__38344;
    wire N__38343;
    wire N__38340;
    wire N__38335;
    wire N__38334;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38317;
    wire N__38312;
    wire N__38309;
    wire N__38308;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38285;
    wire N__38284;
    wire N__38283;
    wire N__38282;
    wire N__38281;
    wire N__38280;
    wire N__38279;
    wire N__38278;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38267;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38255;
    wire N__38252;
    wire N__38249;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38230;
    wire N__38229;
    wire N__38228;
    wire N__38227;
    wire N__38222;
    wire N__38219;
    wire N__38214;
    wire N__38211;
    wire N__38206;
    wire N__38203;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38185;
    wire N__38180;
    wire N__38171;
    wire N__38168;
    wire N__38165;
    wire N__38164;
    wire N__38161;
    wire N__38160;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38148;
    wire N__38141;
    wire N__38138;
    wire N__38135;
    wire N__38132;
    wire N__38129;
    wire N__38128;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38117;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38103;
    wire N__38102;
    wire N__38101;
    wire N__38098;
    wire N__38093;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38069;
    wire N__38066;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38042;
    wire N__38039;
    wire N__38036;
    wire N__38031;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38008;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37997;
    wire N__37996;
    wire N__37993;
    wire N__37990;
    wire N__37987;
    wire N__37984;
    wire N__37983;
    wire N__37980;
    wire N__37979;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37961;
    wire N__37956;
    wire N__37943;
    wire N__37940;
    wire N__37939;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37913;
    wire N__37910;
    wire N__37907;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37892;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37880;
    wire N__37879;
    wire N__37878;
    wire N__37875;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37861;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37853;
    wire N__37852;
    wire N__37847;
    wire N__37844;
    wire N__37841;
    wire N__37838;
    wire N__37835;
    wire N__37832;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37809;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37782;
    wire N__37779;
    wire N__37772;
    wire N__37769;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37759;
    wire N__37756;
    wire N__37753;
    wire N__37752;
    wire N__37751;
    wire N__37746;
    wire N__37743;
    wire N__37740;
    wire N__37739;
    wire N__37736;
    wire N__37735;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37706;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37694;
    wire N__37689;
    wire N__37686;
    wire N__37679;
    wire N__37676;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37658;
    wire N__37655;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37649;
    wire N__37646;
    wire N__37643;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37633;
    wire N__37632;
    wire N__37629;
    wire N__37628;
    wire N__37625;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37615;
    wire N__37612;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37571;
    wire N__37568;
    wire N__37563;
    wire N__37560;
    wire N__37551;
    wire N__37548;
    wire N__37543;
    wire N__37540;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37523;
    wire N__37522;
    wire N__37521;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37490;
    wire N__37487;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37475;
    wire N__37472;
    wire N__37467;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37451;
    wire N__37448;
    wire N__37445;
    wire N__37440;
    wire N__37435;
    wire N__37432;
    wire N__37427;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37406;
    wire N__37403;
    wire N__37400;
    wire N__37397;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37389;
    wire N__37388;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37375;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37352;
    wire N__37351;
    wire N__37344;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37332;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37210;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37184;
    wire N__37181;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37154;
    wire N__37151;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37121;
    wire N__37118;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37108;
    wire N__37105;
    wire N__37100;
    wire N__37097;
    wire N__37096;
    wire N__37095;
    wire N__37094;
    wire N__37093;
    wire N__37092;
    wire N__37091;
    wire N__37090;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37086;
    wire N__37085;
    wire N__37084;
    wire N__37083;
    wire N__37082;
    wire N__37073;
    wire N__37064;
    wire N__37055;
    wire N__37046;
    wire N__37045;
    wire N__37036;
    wire N__37033;
    wire N__37028;
    wire N__37025;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36992;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36984;
    wire N__36979;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36965;
    wire N__36964;
    wire N__36963;
    wire N__36962;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36953;
    wire N__36952;
    wire N__36951;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36943;
    wire N__36940;
    wire N__36939;
    wire N__36938;
    wire N__36937;
    wire N__36936;
    wire N__36935;
    wire N__36934;
    wire N__36933;
    wire N__36930;
    wire N__36929;
    wire N__36928;
    wire N__36927;
    wire N__36922;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36906;
    wire N__36903;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36875;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36851;
    wire N__36846;
    wire N__36845;
    wire N__36844;
    wire N__36843;
    wire N__36842;
    wire N__36841;
    wire N__36840;
    wire N__36839;
    wire N__36838;
    wire N__36837;
    wire N__36836;
    wire N__36835;
    wire N__36834;
    wire N__36833;
    wire N__36832;
    wire N__36831;
    wire N__36830;
    wire N__36829;
    wire N__36828;
    wire N__36827;
    wire N__36826;
    wire N__36825;
    wire N__36824;
    wire N__36823;
    wire N__36822;
    wire N__36821;
    wire N__36820;
    wire N__36819;
    wire N__36818;
    wire N__36817;
    wire N__36816;
    wire N__36815;
    wire N__36814;
    wire N__36813;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36609;
    wire N__36604;
    wire N__36599;
    wire N__36596;
    wire N__36593;
    wire N__36592;
    wire N__36591;
    wire N__36588;
    wire N__36583;
    wire N__36580;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36568;
    wire N__36567;
    wire N__36566;
    wire N__36565;
    wire N__36564;
    wire N__36563;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36553;
    wire N__36552;
    wire N__36551;
    wire N__36550;
    wire N__36547;
    wire N__36546;
    wire N__36545;
    wire N__36544;
    wire N__36543;
    wire N__36540;
    wire N__36539;
    wire N__36532;
    wire N__36527;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36506;
    wire N__36503;
    wire N__36502;
    wire N__36499;
    wire N__36498;
    wire N__36495;
    wire N__36494;
    wire N__36491;
    wire N__36486;
    wire N__36483;
    wire N__36474;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36457;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36439;
    wire N__36422;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36414;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36301;
    wire N__36298;
    wire N__36295;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36272;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36166;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36134;
    wire N__36131;
    wire N__36130;
    wire N__36127;
    wire N__36126;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36114;
    wire N__36111;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36097;
    wire N__36094;
    wire N__36091;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36072;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36055;
    wire N__36054;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36042;
    wire N__36035;
    wire N__36034;
    wire N__36033;
    wire N__36032;
    wire N__36029;
    wire N__36024;
    wire N__36021;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36007;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35984;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35972;
    wire N__35971;
    wire N__35966;
    wire N__35965;
    wire N__35964;
    wire N__35963;
    wire N__35962;
    wire N__35961;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35909;
    wire N__35906;
    wire N__35905;
    wire N__35904;
    wire N__35901;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35885;
    wire N__35882;
    wire N__35879;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35864;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35816;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35809;
    wire N__35808;
    wire N__35807;
    wire N__35806;
    wire N__35805;
    wire N__35796;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35772;
    wire N__35767;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35729;
    wire N__35726;
    wire N__35723;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35696;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35669;
    wire N__35666;
    wire N__35663;
    wire N__35660;
    wire N__35657;
    wire N__35656;
    wire N__35655;
    wire N__35654;
    wire N__35653;
    wire N__35652;
    wire N__35649;
    wire N__35638;
    wire N__35633;
    wire N__35630;
    wire N__35629;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35621;
    wire N__35620;
    wire N__35617;
    wire N__35612;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35585;
    wire N__35582;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35480;
    wire N__35477;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35469;
    wire N__35464;
    wire N__35461;
    wire N__35460;
    wire N__35459;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35426;
    wire N__35425;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35417;
    wire N__35414;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35365;
    wire N__35364;
    wire N__35363;
    wire N__35360;
    wire N__35355;
    wire N__35352;
    wire N__35345;
    wire N__35344;
    wire N__35343;
    wire N__35342;
    wire N__35337;
    wire N__35336;
    wire N__35331;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35303;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35287;
    wire N__35276;
    wire N__35273;
    wire N__35272;
    wire N__35271;
    wire N__35268;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35257;
    wire N__35254;
    wire N__35253;
    wire N__35252;
    wire N__35251;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35236;
    wire N__35231;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35189;
    wire N__35186;
    wire N__35185;
    wire N__35184;
    wire N__35183;
    wire N__35182;
    wire N__35181;
    wire N__35180;
    wire N__35177;
    wire N__35174;
    wire N__35169;
    wire N__35164;
    wire N__35161;
    wire N__35150;
    wire N__35147;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35132;
    wire N__35131;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35120;
    wire N__35117;
    wire N__35112;
    wire N__35109;
    wire N__35102;
    wire N__35099;
    wire N__35098;
    wire N__35097;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35017;
    wire N__35014;
    wire N__35009;
    wire N__35006;
    wire N__35001;
    wire N__34994;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34986;
    wire N__34985;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34975;
    wire N__34974;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34959;
    wire N__34954;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34930;
    wire N__34927;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34916;
    wire N__34913;
    wire N__34908;
    wire N__34907;
    wire N__34904;
    wire N__34903;
    wire N__34898;
    wire N__34895;
    wire N__34894;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34872;
    wire N__34869;
    wire N__34862;
    wire N__34859;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34837;
    wire N__34836;
    wire N__34835;
    wire N__34834;
    wire N__34833;
    wire N__34832;
    wire N__34831;
    wire N__34830;
    wire N__34829;
    wire N__34828;
    wire N__34827;
    wire N__34824;
    wire N__34819;
    wire N__34814;
    wire N__34805;
    wire N__34800;
    wire N__34797;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34753;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34745;
    wire N__34742;
    wire N__34739;
    wire N__34734;
    wire N__34733;
    wire N__34732;
    wire N__34731;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34725;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34708;
    wire N__34703;
    wire N__34696;
    wire N__34693;
    wire N__34686;
    wire N__34683;
    wire N__34676;
    wire N__34673;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34651;
    wire N__34650;
    wire N__34649;
    wire N__34644;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34623;
    wire N__34622;
    wire N__34617;
    wire N__34614;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34600;
    wire N__34595;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34577;
    wire N__34568;
    wire N__34565;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34499;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34484;
    wire N__34481;
    wire N__34476;
    wire N__34473;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34454;
    wire N__34451;
    wire N__34448;
    wire N__34445;
    wire N__34442;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34428;
    wire N__34427;
    wire N__34426;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34367;
    wire N__34362;
    wire N__34357;
    wire N__34352;
    wire N__34351;
    wire N__34350;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34331;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34312;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34300;
    wire N__34299;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34282;
    wire N__34279;
    wire N__34278;
    wire N__34277;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34245;
    wire N__34244;
    wire N__34241;
    wire N__34238;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34195;
    wire N__34188;
    wire N__34181;
    wire N__34178;
    wire N__34177;
    wire N__34174;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34124;
    wire N__34121;
    wire N__34116;
    wire N__34113;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34094;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34070;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34062;
    wire N__34061;
    wire N__34060;
    wire N__34057;
    wire N__34054;
    wire N__34049;
    wire N__34046;
    wire N__34045;
    wire N__34042;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34019;
    wire N__34018;
    wire N__34017;
    wire N__34016;
    wire N__34013;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34001;
    wire N__33992;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33965;
    wire N__33962;
    wire N__33955;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33930;
    wire N__33929;
    wire N__33928;
    wire N__33927;
    wire N__33926;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33890;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33877;
    wire N__33876;
    wire N__33875;
    wire N__33874;
    wire N__33873;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33851;
    wire N__33848;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33830;
    wire N__33823;
    wire N__33818;
    wire N__33807;
    wire N__33802;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33776;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33763;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33742;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33688;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33646;
    wire N__33641;
    wire N__33640;
    wire N__33637;
    wire N__33636;
    wire N__33635;
    wire N__33632;
    wire N__33625;
    wire N__33620;
    wire N__33617;
    wire N__33616;
    wire N__33615;
    wire N__33614;
    wire N__33613;
    wire N__33612;
    wire N__33611;
    wire N__33610;
    wire N__33609;
    wire N__33608;
    wire N__33607;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33595;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33583;
    wire N__33582;
    wire N__33579;
    wire N__33574;
    wire N__33573;
    wire N__33572;
    wire N__33569;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33550;
    wire N__33547;
    wire N__33546;
    wire N__33545;
    wire N__33540;
    wire N__33537;
    wire N__33536;
    wire N__33533;
    wire N__33532;
    wire N__33529;
    wire N__33524;
    wire N__33517;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33499;
    wire N__33496;
    wire N__33479;
    wire N__33478;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33474;
    wire N__33473;
    wire N__33472;
    wire N__33467;
    wire N__33460;
    wire N__33455;
    wire N__33452;
    wire N__33443;
    wire N__33442;
    wire N__33441;
    wire N__33440;
    wire N__33439;
    wire N__33436;
    wire N__33429;
    wire N__33426;
    wire N__33419;
    wire N__33416;
    wire N__33415;
    wire N__33414;
    wire N__33413;
    wire N__33412;
    wire N__33411;
    wire N__33410;
    wire N__33409;
    wire N__33408;
    wire N__33407;
    wire N__33404;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33385;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33370;
    wire N__33367;
    wire N__33360;
    wire N__33359;
    wire N__33358;
    wire N__33357;
    wire N__33356;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33338;
    wire N__33335;
    wire N__33330;
    wire N__33325;
    wire N__33320;
    wire N__33317;
    wire N__33296;
    wire N__33295;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33289;
    wire N__33284;
    wire N__33279;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33265;
    wire N__33262;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33254;
    wire N__33253;
    wire N__33250;
    wire N__33245;
    wire N__33242;
    wire N__33239;
    wire N__33238;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33222;
    wire N__33219;
    wire N__33212;
    wire N__33209;
    wire N__33206;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33193;
    wire N__33188;
    wire N__33185;
    wire N__33184;
    wire N__33183;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33172;
    wire N__33169;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33149;
    wire N__33146;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33131;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33125;
    wire N__33124;
    wire N__33123;
    wire N__33122;
    wire N__33121;
    wire N__33120;
    wire N__33109;
    wire N__33106;
    wire N__33105;
    wire N__33102;
    wire N__33097;
    wire N__33092;
    wire N__33089;
    wire N__33084;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33078;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33059;
    wire N__33054;
    wire N__33051;
    wire N__33046;
    wire N__33041;
    wire N__33038;
    wire N__33029;
    wire N__33024;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__33001;
    wire N__33000;
    wire N__32997;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32964;
    wire N__32961;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32943;
    wire N__32942;
    wire N__32939;
    wire N__32936;
    wire N__32935;
    wire N__32934;
    wire N__32931;
    wire N__32930;
    wire N__32929;
    wire N__32926;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32909;
    wire N__32906;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32881;
    wire N__32880;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32868;
    wire N__32861;
    wire N__32860;
    wire N__32857;
    wire N__32856;
    wire N__32855;
    wire N__32854;
    wire N__32851;
    wire N__32846;
    wire N__32843;
    wire N__32838;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32802;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32790;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32750;
    wire N__32747;
    wire N__32742;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32701;
    wire N__32698;
    wire N__32695;
    wire N__32694;
    wire N__32693;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32666;
    wire N__32665;
    wire N__32664;
    wire N__32663;
    wire N__32660;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32627;
    wire N__32620;
    wire N__32617;
    wire N__32612;
    wire N__32603;
    wire N__32600;
    wire N__32595;
    wire N__32588;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32557;
    wire N__32556;
    wire N__32555;
    wire N__32550;
    wire N__32547;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32536;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32474;
    wire N__32471;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32447;
    wire N__32440;
    wire N__32437;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32419;
    wire N__32414;
    wire N__32411;
    wire N__32406;
    wire N__32403;
    wire N__32396;
    wire N__32393;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32375;
    wire N__32374;
    wire N__32373;
    wire N__32372;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32335;
    wire N__32332;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32313;
    wire N__32308;
    wire N__32305;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32290;
    wire N__32287;
    wire N__32286;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32218;
    wire N__32217;
    wire N__32214;
    wire N__32213;
    wire N__32210;
    wire N__32209;
    wire N__32206;
    wire N__32205;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32147;
    wire N__32140;
    wire N__32135;
    wire N__32126;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32107;
    wire N__32104;
    wire N__32103;
    wire N__32102;
    wire N__32099;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32072;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32048;
    wire N__32045;
    wire N__32036;
    wire N__32033;
    wire N__32032;
    wire N__32031;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32018;
    wire N__32017;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__32000;
    wire N__31997;
    wire N__31996;
    wire N__31991;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31930;
    wire N__31919;
    wire N__31918;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31898;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31873;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31850;
    wire N__31847;
    wire N__31838;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31825;
    wire N__31822;
    wire N__31819;
    wire N__31816;
    wire N__31813;
    wire N__31808;
    wire N__31807;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31784;
    wire N__31783;
    wire N__31782;
    wire N__31781;
    wire N__31778;
    wire N__31771;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31753;
    wire N__31752;
    wire N__31751;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31739;
    wire N__31738;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31732;
    wire N__31727;
    wire N__31722;
    wire N__31721;
    wire N__31720;
    wire N__31719;
    wire N__31718;
    wire N__31711;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31693;
    wire N__31682;
    wire N__31679;
    wire N__31678;
    wire N__31677;
    wire N__31676;
    wire N__31675;
    wire N__31672;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31666;
    wire N__31665;
    wire N__31664;
    wire N__31663;
    wire N__31662;
    wire N__31661;
    wire N__31660;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31631;
    wire N__31624;
    wire N__31619;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31594;
    wire N__31593;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31577;
    wire N__31574;
    wire N__31573;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31556;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31541;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31529;
    wire N__31528;
    wire N__31527;
    wire N__31526;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31522;
    wire N__31519;
    wire N__31514;
    wire N__31511;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31499;
    wire N__31498;
    wire N__31497;
    wire N__31496;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31426;
    wire N__31423;
    wire N__31422;
    wire N__31421;
    wire N__31416;
    wire N__31413;
    wire N__31412;
    wire N__31411;
    wire N__31410;
    wire N__31409;
    wire N__31408;
    wire N__31407;
    wire N__31406;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31396;
    wire N__31391;
    wire N__31386;
    wire N__31381;
    wire N__31378;
    wire N__31373;
    wire N__31370;
    wire N__31365;
    wire N__31362;
    wire N__31355;
    wire N__31354;
    wire N__31353;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31316;
    wire N__31311;
    wire N__31308;
    wire N__31295;
    wire N__31294;
    wire N__31293;
    wire N__31290;
    wire N__31289;
    wire N__31288;
    wire N__31287;
    wire N__31286;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31274;
    wire N__31273;
    wire N__31272;
    wire N__31269;
    wire N__31264;
    wire N__31261;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31238;
    wire N__31235;
    wire N__31230;
    wire N__31227;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31217;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31169;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31145;
    wire N__31142;
    wire N__31139;
    wire N__31136;
    wire N__31133;
    wire N__31130;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31103;
    wire N__31100;
    wire N__31097;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31069;
    wire N__31066;
    wire N__31065;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31053;
    wire N__31050;
    wire N__31043;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31019;
    wire N__31018;
    wire N__31017;
    wire N__31016;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31012;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30992;
    wire N__30991;
    wire N__30990;
    wire N__30989;
    wire N__30988;
    wire N__30987;
    wire N__30986;
    wire N__30985;
    wire N__30984;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30972;
    wire N__30967;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30946;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30932;
    wire N__30929;
    wire N__30926;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30901;
    wire N__30900;
    wire N__30899;
    wire N__30896;
    wire N__30895;
    wire N__30894;
    wire N__30891;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30870;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30852;
    wire N__30849;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30818;
    wire N__30817;
    wire N__30816;
    wire N__30815;
    wire N__30814;
    wire N__30809;
    wire N__30802;
    wire N__30801;
    wire N__30800;
    wire N__30799;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30782;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30752;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30722;
    wire N__30719;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30656;
    wire N__30653;
    wire N__30650;
    wire N__30647;
    wire N__30644;
    wire N__30641;
    wire N__30638;
    wire N__30635;
    wire N__30632;
    wire N__30629;
    wire N__30626;
    wire N__30623;
    wire N__30620;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30602;
    wire N__30599;
    wire N__30596;
    wire N__30593;
    wire N__30590;
    wire N__30587;
    wire N__30584;
    wire N__30583;
    wire N__30582;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30572;
    wire N__30569;
    wire N__30566;
    wire N__30565;
    wire N__30564;
    wire N__30563;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30559;
    wire N__30558;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30538;
    wire N__30531;
    wire N__30524;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30502;
    wire N__30501;
    wire N__30500;
    wire N__30499;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30488;
    wire N__30487;
    wire N__30486;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30449;
    wire N__30444;
    wire N__30439;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30417;
    wire N__30414;
    wire N__30413;
    wire N__30412;
    wire N__30409;
    wire N__30404;
    wire N__30403;
    wire N__30400;
    wire N__30399;
    wire N__30398;
    wire N__30397;
    wire N__30394;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30378;
    wire N__30371;
    wire N__30366;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30302;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30284;
    wire N__30283;
    wire N__30282;
    wire N__30281;
    wire N__30280;
    wire N__30279;
    wire N__30278;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30261;
    wire N__30254;
    wire N__30249;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30223;
    wire N__30222;
    wire N__30221;
    wire N__30220;
    wire N__30219;
    wire N__30214;
    wire N__30211;
    wire N__30204;
    wire N__30197;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30155;
    wire N__30152;
    wire N__30149;
    wire N__30146;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30053;
    wire N__30050;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30011;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29960;
    wire N__29957;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29942;
    wire N__29939;
    wire N__29936;
    wire N__29933;
    wire N__29930;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29867;
    wire N__29864;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29848;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29833;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29810;
    wire N__29809;
    wire N__29806;
    wire N__29803;
    wire N__29798;
    wire N__29795;
    wire N__29792;
    wire N__29791;
    wire N__29790;
    wire N__29789;
    wire N__29788;
    wire N__29787;
    wire N__29786;
    wire N__29785;
    wire N__29784;
    wire N__29783;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29773;
    wire N__29772;
    wire N__29771;
    wire N__29770;
    wire N__29767;
    wire N__29766;
    wire N__29759;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29743;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29726;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29707;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29687;
    wire N__29678;
    wire N__29673;
    wire N__29664;
    wire N__29661;
    wire N__29654;
    wire N__29651;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29636;
    wire N__29633;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29618;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29607;
    wire N__29602;
    wire N__29599;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29576;
    wire N__29575;
    wire N__29574;
    wire N__29573;
    wire N__29572;
    wire N__29571;
    wire N__29570;
    wire N__29569;
    wire N__29566;
    wire N__29563;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29555;
    wire N__29552;
    wire N__29551;
    wire N__29550;
    wire N__29547;
    wire N__29546;
    wire N__29543;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29531;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29516;
    wire N__29515;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29494;
    wire N__29491;
    wire N__29486;
    wire N__29483;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29454;
    wire N__29449;
    wire N__29448;
    wire N__29445;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29402;
    wire N__29401;
    wire N__29396;
    wire N__29393;
    wire N__29390;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29373;
    wire N__29366;
    wire N__29357;
    wire N__29354;
    wire N__29353;
    wire N__29352;
    wire N__29351;
    wire N__29350;
    wire N__29349;
    wire N__29348;
    wire N__29345;
    wire N__29342;
    wire N__29341;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29296;
    wire N__29293;
    wire N__29290;
    wire N__29289;
    wire N__29288;
    wire N__29287;
    wire N__29286;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29268;
    wire N__29265;
    wire N__29260;
    wire N__29255;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29237;
    wire N__29232;
    wire N__29229;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29196;
    wire N__29193;
    wire N__29192;
    wire N__29187;
    wire N__29180;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29157;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29143;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29117;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29105;
    wire N__29102;
    wire N__29101;
    wire N__29100;
    wire N__29099;
    wire N__29098;
    wire N__29095;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29057;
    wire N__29054;
    wire N__29051;
    wire N__29048;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29028;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28959;
    wire N__28954;
    wire N__28947;
    wire N__28944;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28925;
    wire N__28916;
    wire N__28913;
    wire N__28912;
    wire N__28911;
    wire N__28908;
    wire N__28907;
    wire N__28904;
    wire N__28903;
    wire N__28902;
    wire N__28901;
    wire N__28900;
    wire N__28899;
    wire N__28898;
    wire N__28895;
    wire N__28894;
    wire N__28891;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28871;
    wire N__28870;
    wire N__28869;
    wire N__28868;
    wire N__28865;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28838;
    wire N__28835;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28799;
    wire N__28792;
    wire N__28789;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28772;
    wire N__28767;
    wire N__28764;
    wire N__28757;
    wire N__28752;
    wire N__28745;
    wire N__28742;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28694;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28676;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28658;
    wire N__28655;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28621;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28597;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28570;
    wire N__28569;
    wire N__28568;
    wire N__28567;
    wire N__28564;
    wire N__28557;
    wire N__28554;
    wire N__28547;
    wire N__28538;
    wire N__28535;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28517;
    wire N__28514;
    wire N__28511;
    wire N__28508;
    wire N__28507;
    wire N__28506;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28495;
    wire N__28492;
    wire N__28491;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28470;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28460;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28430;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28418;
    wire N__28415;
    wire N__28414;
    wire N__28409;
    wire N__28406;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28377;
    wire N__28374;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28358;
    wire N__28355;
    wire N__28352;
    wire N__28349;
    wire N__28346;
    wire N__28343;
    wire N__28340;
    wire N__28337;
    wire N__28332;
    wire N__28327;
    wire N__28324;
    wire N__28319;
    wire N__28314;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28274;
    wire N__28271;
    wire N__28270;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28244;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28236;
    wire N__28235;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28211;
    wire N__28208;
    wire N__28207;
    wire N__28204;
    wire N__28203;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28184;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28151;
    wire N__28148;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28129;
    wire N__28126;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28114;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28082;
    wire N__28079;
    wire N__28074;
    wire N__28073;
    wire N__28066;
    wire N__28063;
    wire N__28058;
    wire N__28055;
    wire N__28054;
    wire N__28053;
    wire N__28052;
    wire N__28051;
    wire N__28050;
    wire N__28049;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28041;
    wire N__28038;
    wire N__28037;
    wire N__28036;
    wire N__28033;
    wire N__28032;
    wire N__28031;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28006;
    wire N__28005;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27898;
    wire N__27893;
    wire N__27890;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27860;
    wire N__27859;
    wire N__27854;
    wire N__27851;
    wire N__27844;
    wire N__27839;
    wire N__27836;
    wire N__27833;
    wire N__27830;
    wire N__27827;
    wire N__27822;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27785;
    wire N__27784;
    wire N__27779;
    wire N__27776;
    wire N__27775;
    wire N__27774;
    wire N__27773;
    wire N__27772;
    wire N__27771;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27763;
    wire N__27762;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27743;
    wire N__27742;
    wire N__27739;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27652;
    wire N__27647;
    wire N__27644;
    wire N__27641;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27619;
    wire N__27616;
    wire N__27609;
    wire N__27606;
    wire N__27601;
    wire N__27600;
    wire N__27597;
    wire N__27592;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27576;
    wire N__27569;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27541;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27533;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27521;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27497;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27476;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27464;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27434;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27410;
    wire N__27407;
    wire N__27402;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27377;
    wire N__27372;
    wire N__27371;
    wire N__27364;
    wire N__27357;
    wire N__27354;
    wire N__27347;
    wire N__27344;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27320;
    wire N__27319;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27313;
    wire N__27312;
    wire N__27309;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27282;
    wire N__27281;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27230;
    wire N__27227;
    wire N__27222;
    wire N__27217;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27197;
    wire N__27194;
    wire N__27191;
    wire N__27188;
    wire N__27183;
    wire N__27182;
    wire N__27175;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27152;
    wire N__27147;
    wire N__27140;
    wire N__27137;
    wire N__27136;
    wire N__27135;
    wire N__27134;
    wire N__27131;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27106;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27083;
    wire N__27080;
    wire N__27079;
    wire N__27076;
    wire N__27075;
    wire N__27074;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27066;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27033;
    wire N__27030;
    wire N__27025;
    wire N__27022;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26964;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26946;
    wire N__26943;
    wire N__26936;
    wire N__26929;
    wire N__26928;
    wire N__26923;
    wire N__26920;
    wire N__26915;
    wire N__26912;
    wire N__26903;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26882;
    wire N__26881;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26839;
    wire N__26838;
    wire N__26835;
    wire N__26830;
    wire N__26825;
    wire N__26822;
    wire N__26821;
    wire N__26820;
    wire N__26817;
    wire N__26812;
    wire N__26807;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26792;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26761;
    wire N__26760;
    wire N__26759;
    wire N__26758;
    wire N__26757;
    wire N__26756;
    wire N__26755;
    wire N__26754;
    wire N__26753;
    wire N__26752;
    wire N__26751;
    wire N__26750;
    wire N__26741;
    wire N__26730;
    wire N__26721;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26704;
    wire N__26703;
    wire N__26700;
    wire N__26695;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26669;
    wire N__26668;
    wire N__26667;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26648;
    wire N__26645;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26615;
    wire N__26612;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26585;
    wire N__26582;
    wire N__26579;
    wire N__26576;
    wire N__26573;
    wire N__26570;
    wire N__26567;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26536;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26507;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26481;
    wire N__26480;
    wire N__26475;
    wire N__26470;
    wire N__26469;
    wire N__26468;
    wire N__26463;
    wire N__26462;
    wire N__26461;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26444;
    wire N__26439;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26369;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26324;
    wire N__26321;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26297;
    wire N__26296;
    wire N__26295;
    wire N__26294;
    wire N__26291;
    wire N__26290;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26279;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26220;
    wire N__26219;
    wire N__26216;
    wire N__26213;
    wire N__26210;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26189;
    wire N__26186;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26168;
    wire N__26165;
    wire N__26162;
    wire N__26159;
    wire N__26156;
    wire N__26153;
    wire N__26148;
    wire N__26141;
    wire N__26138;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26113;
    wire N__26106;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26090;
    wire N__26085;
    wire N__26080;
    wire N__26071;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26014;
    wire N__26013;
    wire N__26010;
    wire N__26005;
    wire N__26000;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25975;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25963;
    wire N__25960;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25948;
    wire N__25943;
    wire N__25942;
    wire N__25941;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25933;
    wire N__25930;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25903;
    wire N__25900;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25883;
    wire N__25882;
    wire N__25879;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25838;
    wire N__25835;
    wire N__25834;
    wire N__25833;
    wire N__25830;
    wire N__25825;
    wire N__25820;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25801;
    wire N__25800;
    wire N__25799;
    wire N__25798;
    wire N__25797;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25788;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25778;
    wire N__25777;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25766;
    wire N__25765;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25737;
    wire N__25736;
    wire N__25733;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25719;
    wire N__25718;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25701;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25685;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25681;
    wire N__25680;
    wire N__25679;
    wire N__25678;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25661;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25640;
    wire N__25629;
    wire N__25626;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25602;
    wire N__25601;
    wire N__25600;
    wire N__25599;
    wire N__25594;
    wire N__25589;
    wire N__25586;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25580;
    wire N__25575;
    wire N__25570;
    wire N__25567;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25544;
    wire N__25543;
    wire N__25538;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25516;
    wire N__25515;
    wire N__25510;
    wire N__25507;
    wire N__25504;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25487;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25462;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25420;
    wire N__25415;
    wire N__25406;
    wire N__25405;
    wire N__25404;
    wire N__25403;
    wire N__25402;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25396;
    wire N__25391;
    wire N__25382;
    wire N__25379;
    wire N__25378;
    wire N__25375;
    wire N__25374;
    wire N__25371;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25363;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25332;
    wire N__25321;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25300;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25292;
    wire N__25291;
    wire N__25288;
    wire N__25285;
    wire N__25278;
    wire N__25275;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25246;
    wire N__25243;
    wire N__25236;
    wire N__25233;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25216;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25210;
    wire N__25209;
    wire N__25206;
    wire N__25201;
    wire N__25200;
    wire N__25199;
    wire N__25198;
    wire N__25195;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25149;
    wire N__25142;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25045;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25025;
    wire N__25022;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24928;
    wire N__24927;
    wire N__24924;
    wire N__24919;
    wire N__24916;
    wire N__24915;
    wire N__24914;
    wire N__24913;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24901;
    wire N__24896;
    wire N__24891;
    wire N__24884;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24866;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24815;
    wire N__24814;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24802;
    wire N__24801;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24771;
    wire N__24770;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24739;
    wire N__24738;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24614;
    wire N__24609;
    wire N__24604;
    wire N__24597;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24575;
    wire N__24574;
    wire N__24573;
    wire N__24572;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24558;
    wire N__24555;
    wire N__24548;
    wire N__24545;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24537;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24526;
    wire N__24525;
    wire N__24522;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24510;
    wire N__24507;
    wire N__24506;
    wire N__24503;
    wire N__24502;
    wire N__24501;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24483;
    wire N__24482;
    wire N__24481;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24466;
    wire N__24463;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24367;
    wire N__24362;
    wire N__24359;
    wire N__24352;
    wire N__24349;
    wire N__24344;
    wire N__24337;
    wire N__24332;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24307;
    wire N__24306;
    wire N__24305;
    wire N__24304;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24292;
    wire N__24287;
    wire N__24282;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24254;
    wire N__24253;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24245;
    wire N__24244;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24209;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24131;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24022;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__24001;
    wire N__24000;
    wire N__23999;
    wire N__23998;
    wire N__23997;
    wire N__23996;
    wire N__23995;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23991;
    wire N__23990;
    wire N__23989;
    wire N__23988;
    wire N__23987;
    wire N__23984;
    wire N__23983;
    wire N__23982;
    wire N__23981;
    wire N__23980;
    wire N__23979;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23972;
    wire N__23971;
    wire N__23968;
    wire N__23959;
    wire N__23956;
    wire N__23955;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23924;
    wire N__23913;
    wire N__23904;
    wire N__23899;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23887;
    wire N__23886;
    wire N__23885;
    wire N__23884;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23860;
    wire N__23855;
    wire N__23850;
    wire N__23849;
    wire N__23846;
    wire N__23839;
    wire N__23832;
    wire N__23827;
    wire N__23824;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23798;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23764;
    wire N__23763;
    wire N__23760;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23740;
    wire N__23737;
    wire N__23734;
    wire N__23723;
    wire N__23722;
    wire N__23721;
    wire N__23720;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23705;
    wire N__23704;
    wire N__23699;
    wire N__23694;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23672;
    wire N__23671;
    wire N__23668;
    wire N__23667;
    wire N__23664;
    wire N__23663;
    wire N__23662;
    wire N__23659;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23634;
    wire N__23631;
    wire N__23626;
    wire N__23621;
    wire N__23620;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23589;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23495;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23272;
    wire N__23269;
    wire N__23264;
    wire N__23261;
    wire N__23258;
    wire N__23257;
    wire N__23256;
    wire N__23255;
    wire N__23254;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23242;
    wire N__23241;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23210;
    wire N__23209;
    wire N__23208;
    wire N__23207;
    wire N__23204;
    wire N__23201;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23183;
    wire N__23182;
    wire N__23181;
    wire N__23180;
    wire N__23179;
    wire N__23178;
    wire N__23177;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23171;
    wire N__23168;
    wire N__23159;
    wire N__23158;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23143;
    wire N__23142;
    wire N__23141;
    wire N__23140;
    wire N__23139;
    wire N__23138;
    wire N__23133;
    wire N__23130;
    wire N__23123;
    wire N__23114;
    wire N__23107;
    wire N__23096;
    wire N__23095;
    wire N__23094;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23067;
    wire N__23060;
    wire N__23059;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23029;
    wire N__23026;
    wire N__23021;
    wire N__23018;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22993;
    wire N__22990;
    wire N__22989;
    wire N__22988;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22972;
    wire N__22971;
    wire N__22968;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22921;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22809;
    wire N__22806;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22778;
    wire N__22775;
    wire N__22770;
    wire N__22765;
    wire N__22758;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22625;
    wire N__22622;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22588;
    wire N__22585;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22568;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22400;
    wire N__22397;
    wire N__22396;
    wire N__22393;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22361;
    wire N__22358;
    wire N__22357;
    wire N__22356;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22344;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22244;
    wire N__22241;
    wire N__22236;
    wire N__22225;
    wire N__22220;
    wire N__22215;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22199;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22136;
    wire N__22135;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22115;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22097;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22085;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22077;
    wire N__22076;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22032;
    wire N__22029;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__21998;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21986;
    wire N__21981;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21968;
    wire N__21957;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21936;
    wire N__21931;
    wire N__21928;
    wire N__21919;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21898;
    wire N__21897;
    wire N__21894;
    wire N__21889;
    wire N__21886;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21850;
    wire N__21849;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21836;
    wire N__21831;
    wire N__21826;
    wire N__21825;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21812;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21784;
    wire N__21781;
    wire N__21780;
    wire N__21779;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21722;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21695;
    wire N__21690;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21643;
    wire N__21640;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21623;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21613;
    wire N__21612;
    wire N__21609;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21595;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21580;
    wire N__21579;
    wire N__21576;
    wire N__21571;
    wire N__21570;
    wire N__21569;
    wire N__21568;
    wire N__21567;
    wire N__21562;
    wire N__21559;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21543;
    wire N__21538;
    wire N__21535;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21516;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21492;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21476;
    wire N__21473;
    wire N__21468;
    wire N__21465;
    wire N__21460;
    wire N__21457;
    wire N__21454;
    wire N__21449;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21417;
    wire N__21414;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21398;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21376;
    wire N__21375;
    wire N__21374;
    wire N__21373;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21350;
    wire N__21345;
    wire N__21342;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21305;
    wire N__21302;
    wire N__21299;
    wire N__21296;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21278;
    wire N__21275;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21263;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21232;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21214;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21190;
    wire N__21189;
    wire N__21188;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21170;
    wire N__21167;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21135;
    wire N__21130;
    wire N__21127;
    wire N__21116;
    wire N__21115;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21100;
    wire N__21099;
    wire N__21092;
    wire N__21091;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20981;
    wire N__20978;
    wire N__20977;
    wire N__20976;
    wire N__20975;
    wire N__20972;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20948;
    wire N__20941;
    wire N__20938;
    wire N__20935;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20866;
    wire N__20865;
    wire N__20864;
    wire N__20863;
    wire N__20860;
    wire N__20853;
    wire N__20852;
    wire N__20849;
    wire N__20844;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20838;
    wire N__20831;
    wire N__20830;
    wire N__20829;
    wire N__20828;
    wire N__20827;
    wire N__20826;
    wire N__20825;
    wire N__20824;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20806;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20741;
    wire N__20738;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20726;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20640;
    wire N__20639;
    wire N__20638;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20627;
    wire N__20624;
    wire N__20623;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20612;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20522;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20492;
    wire N__20489;
    wire N__20486;
    wire N__20477;
    wire N__20472;
    wire N__20469;
    wire N__20464;
    wire N__20459;
    wire N__20454;
    wire N__20449;
    wire N__20446;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20402;
    wire N__20401;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20393;
    wire N__20390;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20379;
    wire N__20378;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20343;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20315;
    wire N__20314;
    wire N__20309;
    wire N__20306;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20263;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20237;
    wire N__20230;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20211;
    wire N__20206;
    wire N__20203;
    wire N__20198;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20169;
    wire N__20166;
    wire N__20165;
    wire N__20162;
    wire N__20159;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20145;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20131;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20084;
    wire N__20081;
    wire N__20078;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20046;
    wire N__20043;
    wire N__20038;
    wire N__20035;
    wire N__20030;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20014;
    wire N__20005;
    wire N__20002;
    wire N__19997;
    wire N__19994;
    wire N__19991;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19928;
    wire N__19927;
    wire N__19926;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19915;
    wire N__19912;
    wire N__19911;
    wire N__19910;
    wire N__19907;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19665;
    wire N__19662;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19547;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19529;
    wire N__19528;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19504;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19461;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19436;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19386;
    wire N__19385;
    wire N__19384;
    wire N__19383;
    wire N__19382;
    wire N__19381;
    wire N__19380;
    wire N__19379;
    wire N__19378;
    wire N__19377;
    wire N__19376;
    wire N__19375;
    wire N__19374;
    wire N__19373;
    wire N__19372;
    wire N__19371;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19359;
    wire N__19352;
    wire N__19341;
    wire N__19338;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19316;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19302;
    wire N__19301;
    wire N__19300;
    wire N__19299;
    wire N__19298;
    wire N__19297;
    wire N__19296;
    wire N__19291;
    wire N__19284;
    wire N__19279;
    wire N__19276;
    wire N__19267;
    wire N__19266;
    wire N__19253;
    wire N__19250;
    wire N__19241;
    wire N__19238;
    wire N__19229;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19172;
    wire N__19169;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19159;
    wire N__19158;
    wire N__19157;
    wire N__19156;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19140;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19115;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19079;
    wire N__19076;
    wire N__19073;
    wire N__19070;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19046;
    wire N__19043;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__19001;
    wire N__19000;
    wire N__18997;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18980;
    wire N__18979;
    wire N__18978;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18955;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18928;
    wire N__18927;
    wire N__18926;
    wire N__18923;
    wire N__18920;
    wire N__18917;
    wire N__18914;
    wire N__18911;
    wire N__18908;
    wire N__18905;
    wire N__18902;
    wire N__18899;
    wire N__18890;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18886;
    wire N__18885;
    wire N__18882;
    wire N__18877;
    wire N__18874;
    wire N__18869;
    wire N__18860;
    wire N__18859;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18845;
    wire N__18842;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18799;
    wire N__18798;
    wire N__18791;
    wire N__18788;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18752;
    wire N__18749;
    wire N__18748;
    wire N__18747;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18726;
    wire N__18723;
    wire N__18718;
    wire N__18713;
    wire N__18710;
    wire N__18707;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18677;
    wire N__18674;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18647;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18626;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18551;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18517;
    wire N__18514;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18479;
    wire N__18476;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18468;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18452;
    wire N__18451;
    wire N__18446;
    wire N__18445;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18409;
    wire N__18408;
    wire N__18407;
    wire N__18404;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18388;
    wire N__18387;
    wire N__18386;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18353;
    wire N__18350;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18304;
    wire N__18303;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18275;
    wire N__18274;
    wire N__18273;
    wire N__18268;
    wire N__18265;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18240;
    wire N__18237;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18223;
    wire N__18222;
    wire N__18221;
    wire N__18218;
    wire N__18213;
    wire N__18208;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17896;
    wire N__17893;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17849;
    wire N__17846;
    wire N__17843;
    wire N__17840;
    wire N__17837;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17501;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17490;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17479;
    wire N__17476;
    wire N__17475;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17463;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17455;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17443;
    wire N__17440;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17429;
    wire N__17428;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17378;
    wire N__17375;
    wire N__17374;
    wire N__17371;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17355;
    wire N__17352;
    wire N__17351;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17277;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17263;
    wire N__17260;
    wire N__17259;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17215;
    wire N__17214;
    wire N__17211;
    wire N__17206;
    wire N__17203;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17143;
    wire N__17142;
    wire N__17141;
    wire N__17138;
    wire N__17131;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17089;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17072;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17055;
    wire N__17050;
    wire N__17047;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17017;
    wire N__17016;
    wire N__17013;
    wire N__17008;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16966;
    wire N__16965;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16953;
    wire N__16946;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16928;
    wire N__16927;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16904;
    wire N__16901;
    wire N__16900;
    wire N__16897;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16862;
    wire N__16861;
    wire N__16860;
    wire N__16855;
    wire N__16852;
    wire N__16847;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16817;
    wire N__16814;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16565;
    wire N__16562;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16550;
    wire N__16547;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16534;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16400;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16346;
    wire N__16343;
    wire N__16340;
    wire N__16337;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16295;
    wire N__16292;
    wire N__16289;
    wire N__16286;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16262;
    wire N__16259;
    wire N__16256;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16220;
    wire N__16219;
    wire N__16216;
    wire N__16215;
    wire N__16212;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16196;
    wire N__16193;
    wire N__16190;
    wire N__16187;
    wire N__16184;
    wire N__16181;
    wire N__16178;
    wire N__16177;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16165;
    wire N__16164;
    wire N__16161;
    wire N__16160;
    wire N__16159;
    wire N__16158;
    wire N__16157;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16139;
    wire N__16136;
    wire N__16127;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16091;
    wire N__16090;
    wire N__16089;
    wire N__16088;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16073;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16065;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16047;
    wire N__16046;
    wire N__16043;
    wire N__16040;
    wire N__16037;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16012;
    wire N__16009;
    wire N__16008;
    wire N__16007;
    wire N__16006;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15975;
    wire N__15968;
    wire N__15965;
    wire N__15962;
    wire N__15959;
    wire N__15956;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15918;
    wire N__15913;
    wire N__15910;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15893;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15850;
    wire N__15847;
    wire N__15846;
    wire N__15841;
    wire N__15838;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15823;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15682;
    wire N__15677;
    wire N__15672;
    wire N__15669;
    wire N__15664;
    wire N__15661;
    wire N__15654;
    wire N__15647;
    wire N__15644;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15619;
    wire N__15614;
    wire N__15611;
    wire N__15610;
    wire N__15609;
    wire N__15606;
    wire N__15601;
    wire N__15596;
    wire N__15593;
    wire N__15592;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15584;
    wire N__15583;
    wire N__15582;
    wire N__15581;
    wire N__15578;
    wire N__15577;
    wire N__15572;
    wire N__15569;
    wire N__15560;
    wire N__15559;
    wire N__15556;
    wire N__15549;
    wire N__15546;
    wire N__15539;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15531;
    wire N__15530;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15519;
    wire N__15514;
    wire N__15507;
    wire N__15504;
    wire N__15497;
    wire N__15494;
    wire N__15493;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15436;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15425;
    wire N__15424;
    wire N__15423;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15409;
    wire N__15408;
    wire N__15405;
    wire N__15404;
    wire N__15403;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15374;
    wire N__15373;
    wire N__15372;
    wire N__15365;
    wire N__15364;
    wire N__15363;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15312;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15279;
    wire N__15276;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15257;
    wire N__15252;
    wire N__15247;
    wire N__15244;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15122;
    wire N__15119;
    wire N__15116;
    wire N__15113;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14971;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14677;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14609;
    wire N__14608;
    wire N__14607;
    wire N__14606;
    wire N__14605;
    wire N__14604;
    wire N__14599;
    wire N__14590;
    wire N__14585;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14579;
    wire N__14578;
    wire N__14575;
    wire N__14566;
    wire N__14561;
    wire N__14560;
    wire N__14559;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14553;
    wire N__14548;
    wire N__14539;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14531;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14520;
    wire N__14515;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14374;
    wire N__14371;
    wire N__14370;
    wire N__14365;
    wire N__14362;
    wire N__14361;
    wire N__14360;
    wire N__14359;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14351;
    wire N__14350;
    wire N__14349;
    wire N__14346;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14331;
    wire N__14326;
    wire N__14319;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14296;
    wire N__14295;
    wire N__14294;
    wire N__14287;
    wire N__14284;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14276;
    wire N__14275;
    wire N__14274;
    wire N__14273;
    wire N__14272;
    wire N__14269;
    wire N__14264;
    wire N__14257;
    wire N__14252;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14226;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14171;
    wire N__14166;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14149;
    wire N__14146;
    wire N__14141;
    wire N__14140;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14108;
    wire N__14105;
    wire N__14104;
    wire N__14103;
    wire N__14102;
    wire N__14101;
    wire N__14094;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14077;
    wire N__14074;
    wire N__14069;
    wire N__14068;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14036;
    wire N__14033;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14021;
    wire N__14018;
    wire N__14015;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13988;
    wire N__13985;
    wire N__13984;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13973;
    wire N__13972;
    wire N__13969;
    wire N__13968;
    wire N__13961;
    wire N__13960;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13930;
    wire N__13925;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13917;
    wire N__13916;
    wire N__13915;
    wire N__13912;
    wire N__13911;
    wire N__13906;
    wire N__13901;
    wire N__13900;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13873;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13846;
    wire N__13845;
    wire N__13844;
    wire N__13841;
    wire N__13840;
    wire N__13835;
    wire N__13832;
    wire N__13831;
    wire N__13830;
    wire N__13827;
    wire N__13826;
    wire N__13825;
    wire N__13822;
    wire N__13821;
    wire N__13818;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13797;
    wire N__13790;
    wire N__13781;
    wire N__13778;
    wire N__13777;
    wire N__13776;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13768;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13760;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13744;
    wire N__13741;
    wire N__13736;
    wire N__13733;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13701;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13683;
    wire N__13680;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13562;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13552;
    wire N__13549;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13495;
    wire N__13492;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13386;
    wire N__13383;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13360;
    wire N__13359;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13106;
    wire N__13099;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13051;
    wire N__13048;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13038;
    wire N__13037;
    wire N__13030;
    wire N__13027;
    wire N__13022;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12859;
    wire N__12854;
    wire N__12851;
    wire N__12850;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12817;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire VCCG0;
    wire GNDG0;
    wire port_data_rw_0_i;
    wire port_clk_c;
    wire \this_delay_clk.M_pipe_qZ0Z_0 ;
    wire rgb_c_3;
    wire rgb_c_1;
    wire \this_delay_clk.M_pipe_qZ0Z_1 ;
    wire \this_delay_clk.M_pipe_qZ0Z_2 ;
    wire rgb_c_2;
    wire rgb_c_4;
    wire rgb_c_5;
    wire M_this_vga_signals_address_6;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_c3_1 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un82_sum_c3_0_cascade_ ;
    wire M_this_vga_signals_address_1;
    wire \this_vga_signals.SUM_3_1 ;
    wire \this_vga_signals.mult1_un75_sum_axb1 ;
    wire \this_vga_signals.mult1_un82_sum_axbxc3_1_2 ;
    wire \this_vga_signals.un2_hsynclto6_0 ;
    wire \this_vga_signals.un4_hsynclt7_cascade_ ;
    wire \this_vga_signals.hsync_1_1 ;
    wire \this_vga_signals.un4_hsynclt8_0_cascade_ ;
    wire this_vga_signals_hsync_1_i;
    wire this_vga_signals_hvisibility_i;
    wire this_vga_signals_vvisibility_i;
    wire rgb_c_0;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3 ;
    wire \this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ;
    wire M_this_vga_signals_address_2;
    wire \this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_ ;
    wire \this_vga_signals.if_m7_0_o4_1_ns_1 ;
    wire \this_vga_signals.SUM_3_cascade_ ;
    wire \this_vga_signals.mult1_un89_sum_axbxc3_1 ;
    wire \this_vga_signals.mult1_un89_sum_c3_0 ;
    wire M_this_vga_signals_address_0;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ;
    wire \this_vga_signals.mult1_un68_sum_c3_2 ;
    wire \this_vga_signals.mult1_un68_sum_c3_2_cascade_ ;
    wire M_this_vga_signals_address_3;
    wire M_this_vga_signals_address_5;
    wire \this_vga_signals.mult1_un61_sum_axbxc3_2 ;
    wire M_this_vga_signals_address_4;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ;
    wire \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ;
    wire \this_vga_signals.SUM_3 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0 ;
    wire \this_vga_signals.mult1_un54_sum_c3_0_cascade_ ;
    wire \this_vga_signals.if_m1_1 ;
    wire \this_vga_ramdac.N_3139_reto ;
    wire bfn_7_17_0_;
    wire \this_vga_signals.un1_M_hcounter_d_cry_1 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_2 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_3 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_4 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_5 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_6 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_7 ;
    wire \this_vga_signals.un1_M_hcounter_d_cry_8 ;
    wire bfn_7_18_0_;
    wire M_this_oam_ram_read_data_14;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_14 ;
    wire M_this_oam_ram_read_data_15;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_15 ;
    wire \this_ppu.oam_cache.N_823_0 ;
    wire \this_ppu.oam_cache.N_820_0 ;
    wire M_this_oam_ram_read_data_8;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_8 ;
    wire M_this_oam_ram_read_data_9;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_9 ;
    wire M_this_oam_ram_read_data_10;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_10 ;
    wire bfn_7_20_0_;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_0 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_1 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_2 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_3 ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_4 ;
    wire \this_ppu.m71_i_o2_0_cascade_ ;
    wire \this_ppu.m71_i_o2_1 ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_0 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_2 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_1 ;
    wire \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ;
    wire \this_ppu.M_oam_cache_cnt_qZ0Z_3 ;
    wire \this_ppu.oam_cache.N_826_0 ;
    wire \this_ppu.oam_cache.N_824_0 ;
    wire \this_ppu.oam_cache.N_821_0 ;
    wire \this_ppu.oam_cache.N_822_0 ;
    wire \this_ppu.oam_cache.N_819_0 ;
    wire \this_ppu.oam_cache.N_825_0 ;
    wire M_this_oam_ram_read_data_0;
    wire M_this_oam_ram_read_data_6;
    wire M_this_oam_ram_read_data_1;
    wire M_this_oam_ram_read_data_3;
    wire M_this_oam_ram_read_data_7;
    wire M_this_oam_ram_read_data_4;
    wire M_this_oam_ram_read_data_5;
    wire M_this_oam_ram_read_data_2;
    wire \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_ ;
    wire \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4 ;
    wire \this_ppu.m35_i_a2_3_cascade_ ;
    wire \this_ppu.N_802_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_2 ;
    wire \this_vga_signals.un2_hsynclto3_1 ;
    wire \this_vga_signals.un2_hsynclto3_1_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_4 ;
    wire \this_vga_ramdac.M_this_vga_ramdac_en_reto ;
    wire \this_vga_ramdac.i2_mux_cascade_ ;
    wire \this_vga_ramdac.N_3140_reto ;
    wire \this_vga_ramdac.N_24_mux_cascade_ ;
    wire \this_vga_ramdac.N_3138_reto ;
    wire \this_ppu.oam_cache.mem_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_5 ;
    wire \this_vga_signals.M_hcounter_d7lt7_0 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_6 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_8 ;
    wire \this_vga_signals.N_864_cascade_ ;
    wire \this_vga_signals.M_hcounter_qZ0Z_7 ;
    wire \this_vga_ramdac.m16_cascade_ ;
    wire \this_vga_ramdac.N_3141_reto ;
    wire \this_vga_ramdac.m19_cascade_ ;
    wire \this_vga_ramdac.N_3142_reto ;
    wire M_this_vram_read_data_0;
    wire M_this_vram_read_data_2;
    wire M_this_vram_read_data_3;
    wire M_this_vram_read_data_1;
    wire \this_vga_ramdac.m6 ;
    wire \this_ppu.oam_cache.mem_17 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_17 ;
    wire \this_ppu.oam_cache.mem_16 ;
    wire \this_vga_ramdac.i2_mux_0 ;
    wire \this_vga_ramdac.N_3143_reto ;
    wire \this_ppu.oam_cache.mem_18 ;
    wire \this_ppu.N_777_0 ;
    wire \this_ppu.N_776_0 ;
    wire \this_ppu.N_932_0_cascade_ ;
    wire \this_ppu.un1_M_state_q_7_i_0_0_cascade_ ;
    wire \this_ppu.N_775_0 ;
    wire \this_ppu.N_932_0 ;
    wire \this_ppu.N_838_7 ;
    wire \this_ppu.M_this_oam_ram_read_data_i_16 ;
    wire bfn_9_21_0_;
    wire \this_ppu.M_this_oam_ram_read_data_i_17 ;
    wire \this_ppu.un1_oam_data_1_cry_0 ;
    wire \this_ppu.M_this_oam_ram_read_data_i_18 ;
    wire \this_ppu.un1_oam_data_1_cry_1 ;
    wire \this_ppu.m28_e_i_o2_0 ;
    wire \this_ppu.un1_oam_data_1_cry_2 ;
    wire \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_3 ;
    wire \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_4 ;
    wire \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ;
    wire \this_ppu.un1_oam_data_1_cry_5 ;
    wire \this_ppu.un1_oam_data_1_cry_6 ;
    wire \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_21 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_22 ;
    wire M_this_oam_ram_read_data_22;
    wire M_this_oam_ram_read_data_i_22;
    wire M_this_oam_ram_read_data_23;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_23 ;
    wire M_this_oam_ram_read_data_24;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_24 ;
    wire M_this_oam_ram_read_data_25;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_25 ;
    wire M_this_oam_ram_read_data_26;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_26 ;
    wire M_this_oam_ram_write_data_14;
    wire M_this_oam_ram_read_data_30;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_30 ;
    wire M_this_oam_ram_write_data_13;
    wire M_this_oam_ram_write_data_15;
    wire M_this_oam_ram_write_data_18;
    wire M_this_oam_ram_read_data_31;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_31 ;
    wire M_this_oam_ram_write_data_8;
    wire M_this_data_tmp_qZ0Z_3;
    wire M_this_oam_ram_write_data_3;
    wire M_this_oam_ram_read_data_21;
    wire M_this_oam_ram_read_data_i_21;
    wire M_this_data_tmp_qZ0Z_6;
    wire M_this_oam_ram_write_data_6;
    wire M_this_oam_ram_write_data_5;
    wire M_this_oam_ram_write_data_7;
    wire M_this_oam_ram_read_data_28;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_28 ;
    wire M_this_oam_ram_read_data_29;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_29 ;
    wire M_this_oam_ram_write_data_16;
    wire M_this_oam_ram_write_data_22;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_19 ;
    wire M_this_oam_ram_read_data_19;
    wire M_this_oam_ram_read_data_i_19;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_20 ;
    wire M_this_oam_ram_read_data_20;
    wire M_this_oam_ram_read_data_i_20;
    wire M_this_oam_ram_write_data_27;
    wire M_this_oam_ram_write_data_30;
    wire M_this_oam_ram_write_data_17;
    wire M_this_oam_ram_write_data_29;
    wire M_this_oam_ram_write_data_24;
    wire dma_0_i;
    wire \this_ppu.oam_cache.mem_7 ;
    wire \this_ppu.oam_cache.mem_3 ;
    wire \this_ppu.oam_cache.mem_4 ;
    wire this_pixel_clk_M_counter_q_i_1;
    wire this_pixel_clk_M_counter_q_0;
    wire \this_vga_signals.M_hcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_hcounter_qZ0Z_0 ;
    wire N_3_0_cascade_;
    wire \this_vga_signals.M_pcounter_q_i_2_0 ;
    wire \this_vga_signals.M_pcounter_q_3_0 ;
    wire \this_vga_signals.N_1188_1 ;
    wire \this_vga_signals.N_1188_1_cascade_ ;
    wire \this_vga_signals.N_933_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_pcounter_qZ0Z_0 ;
    wire N_2_0;
    wire M_this_vga_signals_pixel_clk_0_0;
    wire N_2_0_cascade_;
    wire N_3_0;
    wire G_462;
    wire \this_ppu.M_oam_cache_read_data_i_16 ;
    wire bfn_10_19_0_;
    wire \this_ppu.M_oam_cache_read_data_i_17 ;
    wire M_this_ppu_spr_addr_4;
    wire \this_ppu.offset_y_cry_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_18 ;
    wire \this_ppu.offset_y_cry_1 ;
    wire M_this_ppu_spr_addr_5;
    wire \this_ppu.oam_cache.mem_10 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_10 ;
    wire \this_ppu.N_836_cascade_ ;
    wire \this_ppu.oam_cache.mem_9 ;
    wire bfn_10_20_0_;
    wire M_this_warmup_qZ0Z_2;
    wire un1_M_this_warmup_d_cry_1;
    wire M_this_warmup_qZ0Z_3;
    wire un1_M_this_warmup_d_cry_2;
    wire M_this_warmup_qZ0Z_4;
    wire un1_M_this_warmup_d_cry_3;
    wire M_this_warmup_qZ0Z_5;
    wire un1_M_this_warmup_d_cry_4;
    wire M_this_warmup_qZ0Z_6;
    wire un1_M_this_warmup_d_cry_5;
    wire M_this_warmup_qZ0Z_7;
    wire un1_M_this_warmup_d_cry_6;
    wire M_this_warmup_qZ0Z_8;
    wire un1_M_this_warmup_d_cry_7;
    wire un1_M_this_warmup_d_cry_8;
    wire M_this_warmup_qZ0Z_9;
    wire bfn_10_21_0_;
    wire M_this_warmup_qZ0Z_10;
    wire un1_M_this_warmup_d_cry_9;
    wire M_this_warmup_qZ0Z_11;
    wire un1_M_this_warmup_d_cry_10;
    wire M_this_warmup_qZ0Z_12;
    wire un1_M_this_warmup_d_cry_11;
    wire M_this_warmup_qZ0Z_13;
    wire un1_M_this_warmup_d_cry_12;
    wire M_this_warmup_qZ0Z_14;
    wire un1_M_this_warmup_d_cry_13;
    wire M_this_warmup_qZ0Z_15;
    wire un1_M_this_warmup_d_cry_14;
    wire M_this_warmup_qZ0Z_16;
    wire un1_M_this_warmup_d_cry_15;
    wire un1_M_this_warmup_d_cry_16;
    wire M_this_warmup_qZ0Z_17;
    wire bfn_10_22_0_;
    wire M_this_warmup_qZ0Z_18;
    wire un1_M_this_warmup_d_cry_17;
    wire M_this_warmup_qZ0Z_19;
    wire un1_M_this_warmup_d_cry_18;
    wire M_this_warmup_qZ0Z_20;
    wire un1_M_this_warmup_d_cry_19;
    wire M_this_warmup_qZ0Z_21;
    wire un1_M_this_warmup_d_cry_20;
    wire M_this_warmup_qZ0Z_22;
    wire un1_M_this_warmup_d_cry_21;
    wire M_this_warmup_qZ0Z_23;
    wire un1_M_this_warmup_d_cry_22;
    wire M_this_warmup_qZ0Z_24;
    wire un1_M_this_warmup_d_cry_23;
    wire un1_M_this_warmup_d_cry_24;
    wire M_this_warmup_qZ0Z_25;
    wire bfn_10_23_0_;
    wire M_this_warmup_qZ0Z_26;
    wire un1_M_this_warmup_d_cry_25;
    wire M_this_warmup_qZ0Z_27;
    wire un1_M_this_warmup_d_cry_26;
    wire un1_M_this_warmup_d_cry_27;
    wire M_this_warmup_qZ0Z_28;
    wire M_this_data_tmp_qZ0Z_8;
    wire M_this_data_tmp_qZ0Z_14;
    wire M_this_data_tmp_qZ0Z_10;
    wire M_this_oam_ram_write_data_10;
    wire M_this_oam_ram_write_data_12;
    wire M_this_data_tmp_qZ0Z_7;
    wire M_this_data_tmp_qZ0Z_5;
    wire M_this_data_tmp_qZ0Z_22;
    wire M_this_data_tmp_qZ0Z_16;
    wire M_this_oam_ram_write_data_31;
    wire M_this_oam_ram_write_data_21;
    wire M_this_oam_ram_write_data_23;
    wire \this_spr_ram.mem_WE_12 ;
    wire \this_spr_ram.mem_WE_14 ;
    wire \this_ppu.oam_cache.mem_5 ;
    wire \this_spr_ram.mem_WE_0 ;
    wire N_34_i;
    wire \this_ppu.oam_cache.mem_14 ;
    wire \this_ppu.M_oam_curr_qc_0_1_cascade_ ;
    wire \this_ppu.m35_i_a2_4 ;
    wire \this_ppu.N_827_0_cascade_ ;
    wire \this_ppu.un1_M_screen_x_q_c2_cascade_ ;
    wire \this_ppu.un1_M_screen_x_q_c5 ;
    wire \this_ppu.un1_M_screen_x_q_c5_cascade_ ;
    wire M_this_ppu_vram_addr_5;
    wire M_this_ppu_vram_addr_6;
    wire \this_ppu.un1_M_screen_x_q_c2 ;
    wire M_this_ppu_vram_addr_1;
    wire M_this_ppu_vram_addr_0;
    wire M_this_ppu_vram_addr_2;
    wire \this_ppu.N_827_0 ;
    wire \this_ppu.un1_M_screen_x_q_c3_cascade_ ;
    wire M_this_ppu_vram_addr_4;
    wire \this_ppu.N_1210_0 ;
    wire \this_ppu.un1_M_screen_x_q_c3 ;
    wire \this_ppu.oam_cache.mem_13 ;
    wire \this_ppu.oam_cache.mem_12 ;
    wire \this_ppu.m13_0_a2_0_0 ;
    wire \this_ppu.N_844_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_1 ;
    wire M_this_warmup_qZ0Z_1;
    wire M_this_warmup_qZ0Z_0;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_9 ;
    wire \this_ppu.M_oam_cache_read_data_16 ;
    wire M_this_ppu_spr_addr_3;
    wire \this_ppu.M_state_qZ0Z_2 ;
    wire M_this_oam_address_qZ0Z_6;
    wire M_this_oam_address_qZ0Z_7;
    wire M_this_data_tmp_qZ0Z_12;
    wire M_this_data_tmp_qZ0Z_15;
    wire M_this_data_tmp_qZ0Z_13;
    wire M_this_oam_ram_write_data_1;
    wire M_this_data_tmp_qZ0Z_20;
    wire M_this_oam_ram_write_data_20;
    wire M_this_oam_ram_write_data_2;
    wire M_this_data_tmp_qZ0Z_9;
    wire M_this_oam_ram_write_data_9;
    wire M_this_oam_ram_write_data_4;
    wire M_this_data_tmp_qZ0Z_11;
    wire M_this_oam_ram_write_data_11;
    wire M_this_data_tmp_qZ0Z_17;
    wire M_this_data_tmp_qZ0Z_23;
    wire M_this_oam_ram_write_data_19;
    wire M_this_oam_ram_write_data_28;
    wire M_this_oam_ram_write_data_25;
    wire \this_spr_ram.mem_out_bus4_1 ;
    wire \this_spr_ram.mem_out_bus0_1 ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ;
    wire \this_spr_ram.mem_out_bus5_1 ;
    wire \this_spr_ram.mem_out_bus1_1 ;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus7_1 ;
    wire \this_spr_ram.mem_out_bus3_1 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus6_1 ;
    wire \this_spr_ram.mem_out_bus2_1 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ;
    wire \this_spr_ram.mem_out_bus4_3 ;
    wire \this_spr_ram.mem_out_bus0_3 ;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ;
    wire M_this_ppu_vram_addr_3;
    wire \this_vga_signals.N_22_0_cascade_ ;
    wire N_856_i;
    wire \this_spr_ram.mem_out_bus5_3 ;
    wire \this_spr_ram.mem_out_bus1_3 ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_ ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3 ;
    wire M_this_spr_ram_read_data_3_cascade_;
    wire N_25_0_i;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_14 ;
    wire \this_spr_ram.mem_out_bus4_2 ;
    wire \this_spr_ram.mem_out_bus0_2 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_6 ;
    wire \this_ppu.M_state_q_inv_1_cascade_ ;
    wire M_this_map_ram_read_data_6;
    wire \this_ppu.m48_i_a2_0 ;
    wire \this_spr_ram.mem_out_bus5_2 ;
    wire \this_spr_ram.mem_out_bus1_2 ;
    wire \this_spr_ram.mem_out_bus7_2 ;
    wire \this_spr_ram.mem_out_bus3_2 ;
    wire \this_spr_ram.mem_out_bus2_2 ;
    wire \this_spr_ram.mem_out_bus6_2 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_ ;
    wire \this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ;
    wire \this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ;
    wire this_ppu_N_247;
    wire \this_vga_signals.N_22_0 ;
    wire M_this_spr_ram_read_data_2_cascade_;
    wire N_28_0_i;
    wire M_this_ppu_oam_addr_4;
    wire M_this_spr_ram_read_data_2;
    wire M_this_spr_ram_read_data_1;
    wire M_this_spr_ram_read_data_3;
    wire \this_ppu.M_oam_curr_dZ0Z25_cascade_ ;
    wire \this_ppu.N_834_0 ;
    wire M_this_ppu_oam_addr_0;
    wire \this_ppu.N_834_0_cascade_ ;
    wire \this_ppu.un1_M_state_q_7_i_0_0 ;
    wire \this_ppu.un1_M_oam_curr_q_1_c1 ;
    wire M_this_ppu_oam_addr_1;
    wire \this_ppu.un1_M_oam_curr_q_1_c1_cascade_ ;
    wire M_this_ppu_oam_addr_2;
    wire \this_ppu.un1_M_oam_curr_q_1_c3 ;
    wire M_this_ppu_oam_addr_3;
    wire \this_ppu.un1_M_oam_curr_q_1_c3_cascade_ ;
    wire \this_ppu.N_778_0 ;
    wire \this_ppu.un1_M_oam_curr_q_1_c5 ;
    wire M_this_ppu_oam_addr_5;
    wire \this_ppu.M_oam_curr_qc_0_1 ;
    wire \this_ppu.M_oam_curr_qZ0Z_6 ;
    wire M_this_status_flags_qZ0Z_0;
    wire \this_ppu.oam_cache.mem_15 ;
    wire \this_ppu.N_784_0 ;
    wire \this_vga_signals.N_859_cascade_ ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_13 ;
    wire \this_ppu.m9_0_a2_5_cascade_ ;
    wire \this_vga_signals.i22_mux ;
    wire \this_vga_signals.M_lcounter_qZ0Z_1 ;
    wire \this_vga_signals.M_lcounter_qZ0Z_0 ;
    wire \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2 ;
    wire \this_ppu.N_814_cascade_ ;
    wire \this_ppu.N_806_cascade_ ;
    wire \this_ppu.N_806 ;
    wire bfn_12_20_0_;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_0 ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_1 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_3 ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_2 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_4 ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_3 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_5 ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_4 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_6 ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_5 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_6 ;
    wire \this_ppu.M_state_q_RNISP3R6_1Z0Z_10 ;
    wire M_this_oam_ram_read_data_11;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_11 ;
    wire \this_ppu.M_state_q_RNISP3R6Z0Z_10 ;
    wire M_this_oam_address_qZ0Z_3;
    wire M_this_oam_address_qZ0Z_2;
    wire un1_M_this_oam_address_q_c4;
    wire M_this_oam_address_qZ0Z_5;
    wire un1_M_this_oam_address_q_c4_cascade_;
    wire M_this_oam_address_qZ0Z_4;
    wire un1_M_this_oam_address_q_c6;
    wire N_1240_0;
    wire M_this_oam_ram_write_data_0_sqmuxa_cascade_;
    wire M_this_oam_ram_write_data_26;
    wire M_this_oam_ram_write_data_0_sqmuxa;
    wire M_this_oam_ram_write_data_0;
    wire M_this_data_tmp_qZ0Z_0;
    wire M_this_data_tmp_qZ0Z_4;
    wire M_this_data_tmp_qZ0Z_2;
    wire M_this_data_tmp_qZ0Z_21;
    wire \this_spr_ram.mem_out_bus7_0 ;
    wire \this_spr_ram.mem_out_bus3_0 ;
    wire \this_spr_ram.mem_out_bus4_0 ;
    wire \this_spr_ram.mem_out_bus0_0 ;
    wire \this_spr_ram.mem_out_bus5_0 ;
    wire \this_spr_ram.mem_out_bus1_0 ;
    wire \this_spr_ram.mem_out_bus6_0 ;
    wire \this_spr_ram.mem_out_bus2_0 ;
    wire \this_spr_ram.mem_radregZ0Z_12 ;
    wire \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ;
    wire \this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ;
    wire \this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ;
    wire \this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ;
    wire \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ;
    wire M_this_spr_ram_read_data_0;
    wire M_this_map_ram_read_data_7;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_3 ;
    wire M_this_map_ram_read_data_3;
    wire M_this_ppu_spr_addr_9;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_4 ;
    wire M_this_map_ram_read_data_4;
    wire M_this_ppu_spr_addr_10;
    wire M_this_ppu_spr_addr_0;
    wire \this_spr_ram.mem_out_bus6_3 ;
    wire \this_spr_ram.mem_out_bus2_3 ;
    wire \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_5 ;
    wire M_this_map_ram_read_data_5;
    wire \this_spr_ram.mem_radregZ0Z_11 ;
    wire \this_ppu.N_797 ;
    wire \this_ppu.un3_M_screen_y_d_0_c4_cascade_ ;
    wire \this_ppu.N_802 ;
    wire \this_spr_ram.mem_out_bus7_3 ;
    wire \this_spr_ram.mem_out_bus3_3 ;
    wire \this_spr_ram.mem_radregZ0Z_13 ;
    wire \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ;
    wire \this_ppu.M_state_qZ0Z_5 ;
    wire \this_ppu.N_796_0 ;
    wire \this_ppu.M_state_qZ0Z_8 ;
    wire \this_ppu.un1_M_surface_x_q_c6_cascade_ ;
    wire \this_ppu.N_798_0_cascade_ ;
    wire \this_ppu.un1_M_surface_x_q_c3 ;
    wire \this_ppu.un1_M_surface_x_q_c3_cascade_ ;
    wire \this_ppu.N_798_0 ;
    wire \this_ppu.un1_M_surface_x_q_c2_cascade_ ;
    wire \this_ppu.un1_M_surface_x_q_c5_cascade_ ;
    wire \this_ppu.N_800 ;
    wire \this_ppu.N_800_cascade_ ;
    wire \this_ppu.M_state_qZ0Z_11 ;
    wire N_18;
    wire \this_ppu.un1_M_surface_x_q_c2 ;
    wire \this_ppu.M_oam_curr_dZ0Z25 ;
    wire \this_ppu.M_state_qZ0Z_7 ;
    wire \this_ppu.M_state_qZ0Z_9 ;
    wire \this_ppu.un1_M_surface_x_q_c1_cascade_ ;
    wire M_this_scroll_qZ0Z_10;
    wire M_this_scroll_qZ0Z_11;
    wire M_this_scroll_qZ0Z_13;
    wire M_this_scroll_qZ0Z_14;
    wire M_this_scroll_qZ0Z_8;
    wire N_829_0_cascade_;
    wire N_58_0_cascade_;
    wire \this_ppu.N_97_mux ;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_ ;
    wire \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_2 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_1 ;
    wire \this_ppu.M_pixel_cnt_qZ0Z_7 ;
    wire \this_ppu.m9_0_a2_4 ;
    wire \this_ppu.M_pixel_cnt_qZ1Z_0 ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_axb_0 ;
    wire \this_ppu.M_state_q_RNISP3R6_2Z0Z_10 ;
    wire \this_ppu.M_state_q_RNISP3R6_4Z0Z_10 ;
    wire \this_ppu.M_state_q_RNISP3R6_0Z0Z_10 ;
    wire \this_ppu.M_state_qZ0Z_4 ;
    wire \this_ppu.M_state_qZ0Z_10 ;
    wire \this_ppu.N_835_0_cascade_ ;
    wire \this_ppu.N_783_cascade_ ;
    wire \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0 ;
    wire \this_ppu.oam_cache.mem_2 ;
    wire \this_ppu.N_60_0 ;
    wire \this_ppu.M_state_qZ0Z_0 ;
    wire \this_ppu.N_835_0 ;
    wire \this_ppu.N_807 ;
    wire \this_ppu.N_814 ;
    wire \this_ppu.N_783 ;
    wire \this_ppu.M_state_q_RNISP3R6_3Z0Z_10 ;
    wire un1_M_this_oam_address_q_c2;
    wire M_this_data_tmp_qZ0Z_18;
    wire M_this_data_tmp_qZ0Z_1;
    wire M_this_data_tmp_qZ0Z_19;
    wire N_1232_0;
    wire \this_ppu.un3_M_screen_y_d_0_c6 ;
    wire \this_ppu.un3_M_screen_y_d_0_c4 ;
    wire this_ppu_M_screen_y_q_3;
    wire \this_ppu.un3_M_screen_y_d_0_c2 ;
    wire this_ppu_M_screen_y_q_4;
    wire \this_ppu.M_state_qZ0Z_6 ;
    wire \this_ppu.m68_0_a2_2_cascade_ ;
    wire \this_ppu.M_state_q_ns_7 ;
    wire M_this_ppu_vga_is_drawing_cascade_;
    wire this_ppu_M_screen_y_q_5;
    wire this_ppu_M_screen_y_q_6;
    wire \this_ppu.un1_M_surface_x_q_c1 ;
    wire M_this_scroll_qZ0Z_9;
    wire M_this_scroll_qZ0Z_15;
    wire \this_ppu.un1_M_surface_x_q_ac0_11 ;
    wire M_this_scroll_qZ0Z_12;
    wire \this_ppu.un1_M_surface_x_q_c4 ;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_2 ;
    wire M_this_map_ram_read_data_2;
    wire M_this_ppu_spr_addr_8;
    wire bfn_14_18_0_;
    wire \this_ppu.M_screen_y_q_RNICCMV8Z0Z_0 ;
    wire \this_ppu.offset_y ;
    wire \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ;
    wire \this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1 ;
    wire \this_ppu.M_surface_y_qZ0Z_1 ;
    wire \this_ppu.un1_M_surface_y_d_cry_0 ;
    wire \this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2 ;
    wire \this_ppu.M_surface_y_qZ0Z_2 ;
    wire \this_ppu.un1_M_surface_y_d_cry_1 ;
    wire \this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3 ;
    wire M_this_ppu_map_addr_5;
    wire \this_ppu.un1_M_surface_y_d_cry_2 ;
    wire \this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4 ;
    wire M_this_ppu_map_addr_6;
    wire \this_ppu.un1_M_surface_y_d_cry_3 ;
    wire \this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5 ;
    wire M_this_ppu_map_addr_7;
    wire \this_ppu.un1_M_surface_y_d_cry_4 ;
    wire \this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6 ;
    wire M_this_ppu_map_addr_8;
    wire \this_ppu.un1_M_surface_y_d_cry_5 ;
    wire \this_ppu.un1_M_surface_y_d_cry_6 ;
    wire \this_ppu.M_screen_y_qZ0Z_7 ;
    wire bfn_14_19_0_;
    wire M_this_ppu_map_addr_9;
    wire M_this_ppu_vram_addr_7;
    wire \this_ppu.M_screen_y_qZ0Z_1 ;
    wire M_this_ppu_vga_is_drawing;
    wire \this_ppu.M_screen_y_qZ0Z_2 ;
    wire \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0 ;
    wire M_this_oam_ram_read_data_12;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_12 ;
    wire \this_delay_clk.M_pipe_qZ0Z_3 ;
    wire N_1256_0;
    wire M_this_oam_ram_read_data_16;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_16 ;
    wire M_this_oam_ram_read_data_17;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_17 ;
    wire M_this_oam_ram_read_data_18;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_18 ;
    wire M_this_oam_ram_read_data_27;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_27 ;
    wire M_this_ctrl_flags_qZ0Z_6;
    wire M_this_oam_ram_read_data_13;
    wire \this_ppu.M_state_qZ0Z_3 ;
    wire \this_ppu.oam_cache.M_oam_cache_write_data_13 ;
    wire M_this_oam_address_qZ0Z_1;
    wire M_this_oam_address_qZ0Z_0;
    wire N_222_0;
    wire N_1248_0;
    wire \this_reset_cond.M_stage_qZ0Z_2 ;
    wire M_this_spr_ram_write_en_0_i_1_0_cascade_;
    wire \this_spr_ram.mem_WE_2 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0 ;
    wire \this_vga_signals.M_vcounter_d7lt8_0_cascade_ ;
    wire \this_ppu.offset_x ;
    wire \this_ppu.M_oam_cache_read_data_i_8 ;
    wire bfn_15_17_0_;
    wire \this_ppu.M_oam_cache_read_data_i_9 ;
    wire \this_ppu.M_surface_x_qZ0Z_1 ;
    wire M_this_ppu_spr_addr_1;
    wire \this_ppu.offset_x_cry_0 ;
    wire \this_ppu.M_oam_cache_read_data_i_10 ;
    wire \this_ppu.M_surface_x_qZ0Z_2 ;
    wire M_this_ppu_spr_addr_2;
    wire \this_ppu.offset_x_cry_1 ;
    wire M_this_ppu_map_addr_0;
    wire \this_ppu.offset_x_3 ;
    wire \this_ppu.offset_x_cry_2 ;
    wire M_this_ppu_map_addr_1;
    wire \this_ppu.offset_x_4 ;
    wire \this_ppu.offset_x_cry_3 ;
    wire \this_ppu.M_oam_cache_read_data_i_13 ;
    wire M_this_ppu_map_addr_2;
    wire \this_ppu.offset_x_5 ;
    wire \this_ppu.offset_x_cry_4 ;
    wire \this_ppu.M_oam_cache_read_data_i_14 ;
    wire M_this_ppu_map_addr_3;
    wire \this_ppu.offset_x_6 ;
    wire \this_ppu.offset_x_cry_5 ;
    wire M_this_ppu_map_addr_4;
    wire \this_ppu.M_oam_cache_read_data_15 ;
    wire \this_ppu.offset_x_cry_6 ;
    wire \this_ppu.offset_x_7 ;
    wire M_this_scroll_qZ0Z_0;
    wire M_this_scroll_qZ0Z_1;
    wire M_this_scroll_qZ0Z_2;
    wire M_this_scroll_qZ0Z_3;
    wire M_this_scroll_qZ0Z_4;
    wire M_this_scroll_qZ0Z_5;
    wire M_this_scroll_qZ0Z_6;
    wire M_this_scroll_qZ0Z_7;
    wire bfn_15_19_0_;
    wire M_this_data_count_q_cry_0_THRU_CO;
    wire M_this_data_count_q_cry_0;
    wire M_this_data_count_q_cry_1_THRU_CO;
    wire M_this_data_count_q_cry_1;
    wire M_this_data_count_q_cry_2_THRU_CO;
    wire M_this_data_count_q_cry_2;
    wire M_this_data_count_q_cry_3;
    wire M_this_data_count_q_cry_4;
    wire M_this_data_count_q_cry_5;
    wire M_this_data_count_q_cry_6_THRU_CO;
    wire M_this_data_count_q_cry_6;
    wire M_this_data_count_q_cry_7;
    wire bfn_15_20_0_;
    wire M_this_data_count_q_cry_8;
    wire M_this_data_count_q_cry_9;
    wire M_this_data_count_q_cry_10;
    wire CONSTANT_ONE_NET;
    wire M_this_data_count_q_cry_11;
    wire M_this_data_count_q_cry_12;
    wire port_enb_c;
    wire M_this_delay_clk_out_0;
    wire M_this_data_count_q_s_8;
    wire N_92;
    wire M_this_data_count_qZ0Z_8;
    wire M_this_data_count_q_cry_3_THRU_CO;
    wire M_this_data_count_qZ0Z_4;
    wire M_this_data_count_q_cry_4_THRU_CO;
    wire M_this_data_count_qZ0Z_5;
    wire M_this_data_count_q_cry_8_THRU_CO;
    wire M_this_data_count_qZ0Z_9;
    wire \this_start_data_delay.M_last_qZ0 ;
    wire N_685_i_cascade_;
    wire M_this_data_count_qZ0Z_2;
    wire M_this_data_count_qZ0Z_1;
    wire M_this_data_count_qZ0Z_3;
    wire M_this_data_count_qZ0Z_0;
    wire \this_reset_cond.M_stage_qZ0Z_1 ;
    wire \this_reset_cond.M_stage_qZ0Z_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_4 ;
    wire \this_reset_cond.M_stage_qZ0Z_0 ;
    wire M_this_map_ram_read_data_0;
    wire M_this_ppu_spr_addr_6;
    wire \this_ppu.oam_cache.mem_0 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ;
    wire bfn_16_15_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_1 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_2 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7 ;
    wire bfn_16_16_0_;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8 ;
    wire \this_vga_signals.M_vcounter_d7lto9_i_a2_1 ;
    wire port_nmib_1_i;
    wire \this_ppu.M_oam_cache_read_data_i_11 ;
    wire \this_ppu.oam_cache.mem_11 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_11 ;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_12 ;
    wire \this_ppu.M_oam_cache_read_data_i_12 ;
    wire \this_ppu.oam_cache.mem_8 ;
    wire \this_ppu.M_oam_cache_read_data_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_0 ;
    wire \this_vga_signals.N_3_1_cascade_ ;
    wire \this_vga_signals.g0_41_N_2L1 ;
    wire \this_vga_signals.g0_41_N_4L5_cascade_ ;
    wire \this_vga_signals.g0_41_1 ;
    wire M_this_vga_ramdac_en;
    wire \this_vga_signals.mult1_un82_sum_c3_0_0_0_1 ;
    wire M_this_vga_signals_address_7;
    wire \this_vga_signals.M_vcounter_qZ0Z_1 ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_ ;
    wire \this_vga_signals.g0_i_x2_4 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_ ;
    wire \this_vga_signals.N_17_i ;
    wire M_this_data_count_q_s_10;
    wire M_this_data_count_q_cry_11_THRU_CO;
    wire M_this_data_count_q_s_13;
    wire M_this_data_count_q_cry_10_THRU_CO;
    wire M_this_data_count_qZ0Z_7;
    wire \this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11 ;
    wire \this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_ ;
    wire \this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11 ;
    wire M_this_data_count_qZ0Z_12;
    wire M_this_data_count_qZ0Z_11;
    wire M_this_data_count_qZ0Z_13;
    wire M_this_data_count_qZ0Z_10;
    wire \this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11 ;
    wire M_this_data_count_q_cry_5_THRU_CO;
    wire N_685_i;
    wire M_this_data_count_qZ0Z_6;
    wire M_this_ctrl_flags_qZ0Z_5;
    wire M_this_ctrl_flags_qZ0Z_7;
    wire \this_reset_cond.M_stage_qZ0Z_5 ;
    wire M_this_spr_address_qZ0Z_0;
    wire bfn_17_12_0_;
    wire M_this_spr_address_qZ0Z_1;
    wire un1_M_this_spr_address_q_cry_0;
    wire M_this_spr_address_qZ0Z_2;
    wire un1_M_this_spr_address_q_cry_1;
    wire M_this_spr_address_qZ0Z_3;
    wire un1_M_this_spr_address_q_cry_2;
    wire M_this_spr_address_qZ0Z_4;
    wire un1_M_this_spr_address_q_cry_3;
    wire M_this_spr_address_qZ0Z_5;
    wire un1_M_this_spr_address_q_cry_4;
    wire M_this_spr_address_qZ0Z_6;
    wire un1_M_this_spr_address_q_cry_5;
    wire M_this_spr_address_qZ0Z_7;
    wire un1_M_this_spr_address_q_cry_6;
    wire un1_M_this_spr_address_q_cry_7;
    wire M_this_spr_address_qZ0Z_8;
    wire bfn_17_13_0_;
    wire M_this_spr_address_qZ0Z_9;
    wire un1_M_this_spr_address_q_cry_8;
    wire M_this_spr_address_qZ0Z_10;
    wire un1_M_this_spr_address_q_cry_9;
    wire un1_M_this_spr_address_q_cry_10;
    wire un1_M_this_spr_address_q_cry_11;
    wire un1_M_this_spr_address_q_cry_12;
    wire M_this_spr_ram_write_en_0_i_1;
    wire \this_vga_signals.M_vcounter_d8 ;
    wire \this_vga_signals.M_hcounter_d7_0 ;
    wire \this_vga_signals.m43_5 ;
    wire this_vga_signals_vsync_1_i;
    wire N_52_0;
    wire N_58_0;
    wire \this_ppu.line_clk.M_last_qZ0 ;
    wire \this_vga_signals.GZ0Z_424 ;
    wire \this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9 ;
    wire \this_ppu.oam_cache.mem_1 ;
    wire \this_vga_signals.vvisibility_0_cascade_ ;
    wire \this_vga_signals.vvisibility ;
    wire \this_vga_signals.g0_0_i_0_1 ;
    wire \this_vga_signals.N_10_i_cascade_ ;
    wire \this_vga_signals.g2_1_2 ;
    wire \this_vga_signals.N_10_i_0 ;
    wire \this_vga_signals.g0_0_i_0_cascade_ ;
    wire \this_vga_signals.if_m5_i_0_0 ;
    wire \this_vga_signals.mult1_un68_sum_c3_0_0_0 ;
    wire \this_vga_signals.if_N_10_0_0_0 ;
    wire \this_vga_signals.g0_1_0_3 ;
    wire \this_vga_signals.g0_1_1_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ;
    wire \this_vga_signals.g0_41_N_3L3_1 ;
    wire \this_vga_signals.mult1_un54_sum_c3_x0_cascade_ ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_;
    wire \this_vga_signals.g0_41_N_4L5_1 ;
    wire N_6_i;
    wire \this_vga_signals.g0_1_1_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c2_0_0 ;
    wire \this_vga_signals.g1_4 ;
    wire \this_vga_signals.g1_0_0_0 ;
    wire \this_vga_signals.g1_0_1_0_cascade_ ;
    wire \this_vga_signals.N_10 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_2_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_ ;
    wire \this_vga_signals.N_5_i_0_cascade_ ;
    wire \this_vga_signals.g1_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ;
    wire \this_vga_signals.g0_i_x2_1 ;
    wire GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO;
    wire \this_spr_ram.mem_WE_8 ;
    wire \this_vga_signals.m43_4 ;
    wire \this_vga_signals.vaddress_c3_d_0 ;
    wire \this_vga_signals.g0_1_0_1 ;
    wire \this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_ ;
    wire \this_vga_signals.CO0_0_i_i_cascade_ ;
    wire \this_vga_signals.vaddress_c5_a0_0_cascade_ ;
    wire \this_vga_signals.vaddress_9_cascade_ ;
    wire \this_vga_signals.g1_3_0_cascade_ ;
    wire \this_vga_signals.N_5_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_c3_0_0_0 ;
    wire \this_vga_signals.N_4_1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_c3_x1 ;
    wire \this_vga_signals.mult1_un54_sum_c2_0_cascade_ ;
    wire \this_vga_signals.g1_1_0_0_cascade_ ;
    wire \this_vga_signals.N_20_0 ;
    wire \this_vga_signals.g0_2_0_3_cascade_ ;
    wire \this_vga_signals.g0_0_0_1_0 ;
    wire \this_vga_signals.g0_0_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4 ;
    wire \this_vga_signals.g0_2_0_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_4 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0 ;
    wire \this_vga_signals.g0_6_0 ;
    wire \this_vga_signals.g0_0_0_1 ;
    wire \this_vga_signals.g0_5_5_N_2L1 ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0;
    wire \this_vga_signals.g0_5_0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3 ;
    wire \this_vga_signals.g1_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_d_0 ;
    wire \this_vga_signals.g0_1_0_cascade_ ;
    wire \this_vga_signals.N_7_1_0_2 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ;
    wire \this_vga_signals.g3_1 ;
    wire \this_vga_signals.g1_3 ;
    wire \this_vga_signals.N_7_1_0_0 ;
    wire \this_vga_signals.g0_1_0_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_ns ;
    wire \this_vga_signals.g1_0 ;
    wire \this_vga_signals.mult1_un54_sum_c2_0 ;
    wire \this_vga_signals.g0_29_1 ;
    wire \this_vga_signals.g1_0_cascade_ ;
    wire this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0;
    wire \this_vga_signals.g0_3 ;
    wire \this_reset_cond.M_stage_qZ0Z_6 ;
    wire M_this_reset_cond_out_0;
    wire rst_n_c;
    wire \this_reset_cond.M_stage_qZ0Z_7 ;
    wire \this_reset_cond.M_stage_qZ0Z_8 ;
    wire \this_spr_ram.mem_WE_10 ;
    wire \this_vga_signals.N_12_0_0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_4 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_5 ;
    wire \this_vga_signals.vaddress_c2_cascade_ ;
    wire \this_vga_signals.N_7_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0 ;
    wire \this_vga_signals.g0_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_x0 ;
    wire \this_vga_signals.vaddress_ac0_9_0_a0_1 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc1 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_ ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_ ;
    wire \this_vga_signals.g0_5_5 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_3 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_2 ;
    wire \this_vga_signals.N_5_i_1 ;
    wire \this_vga_signals.N_5786_0_0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x0 ;
    wire \this_vga_signals.mult1_un47_sum_axbxc3_x1 ;
    wire \this_vga_signals.CO0_0_i_i ;
    wire \this_vga_signals.N_12_0 ;
    wire \this_vga_signals.N_12_0_cascade_ ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ;
    wire \this_vga_signals.mult1_un61_sum_axb1_0_1 ;
    wire \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_x0 ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_ns ;
    wire \this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_ ;
    wire \this_vga_signals.mult1_un54_sum_axbxc3_1 ;
    wire \this_vga_signals.g0_2_0_1 ;
    wire \this_vga_signals.mult1_un54_sum_axb1_out_0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ;
    wire port_rw_in;
    wire M_this_state_d_0_sqmuxa_2_cascade_;
    wire \this_start_data_delay.N_233_0_cascade_ ;
    wire N_164;
    wire \this_vga_signals.g1_3_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6 ;
    wire \this_spr_ram.mem_WE_6 ;
    wire M_this_spr_address_qZ0Z_12;
    wire M_this_spr_address_qZ0Z_11;
    wire M_this_spr_address_qZ0Z_13;
    wire M_this_spr_ram_write_en_0_i_1_0;
    wire \this_spr_ram.mem_WE_4 ;
    wire M_this_spr_ram_write_data_3;
    wire \this_ppu.oam_cache.M_oam_cache_read_data_1 ;
    wire M_this_map_ram_read_data_1;
    wire \this_ppu.M_state_q_inv_1 ;
    wire M_this_ppu_spr_addr_7;
    wire M_this_spr_ram_write_data_1;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ;
    wire \this_vga_signals.mult1_un40_sum_c3_0 ;
    wire \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_ ;
    wire \this_vga_signals.N_14 ;
    wire \this_vga_signals.g1_6 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_5 ;
    wire \this_vga_signals.N_7_1_0_3_cascade_ ;
    wire \this_vga_signals.G_5_i_o2_0_1 ;
    wire \this_vga_signals.vaddress_8 ;
    wire \this_vga_signals.vaddress_9 ;
    wire \this_vga_signals.N_19_0_0 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_6 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_9 ;
    wire \this_vga_signals.m47_0_0 ;
    wire \this_vga_signals.m47_0_1_cascade_ ;
    wire this_vga_signals_M_vcounter_q_6;
    wire \this_vga_signals.M_vcounter_qZ0Z_4 ;
    wire \this_vga_signals.SUM_2_cascade_ ;
    wire \this_vga_signals.g0_0_i_a7_1 ;
    wire N_88;
    wire port_address_in_5;
    wire port_address_in_7;
    wire port_address_in_3;
    wire \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ;
    wire \this_vga_signals.M_vcounter_q_4_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_5_repZ0Z1 ;
    wire \this_vga_signals.vaddress_7 ;
    wire \this_vga_signals.vaddress_6 ;
    wire \this_vga_signals.vaddress_5 ;
    wire \this_vga_signals.vaddress_7_cascade_ ;
    wire \this_vga_signals.SUM_2 ;
    wire \this_vga_signals.if_m2_0 ;
    wire \this_start_data_delay.N_345_cascade_ ;
    wire \this_start_data_delay.N_284_0 ;
    wire \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_ ;
    wire \this_start_data_delay.N_23_1_0_cascade_ ;
    wire \this_start_data_delay.N_339_cascade_ ;
    wire \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6 ;
    wire M_this_substate_qZ0;
    wire \this_start_data_delay.N_467 ;
    wire \this_start_data_delay.N_386_cascade_ ;
    wire port_address_in_1;
    wire \this_start_data_delay.N_380 ;
    wire \this_start_data_delay.N_341 ;
    wire M_this_spr_ram_write_data_2;
    wire dma_axb0_cascade_;
    wire dma_0;
    wire dma_axb3;
    wire \this_vga_signals.vaddress_c2 ;
    wire \this_vga_signals.N_13 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ;
    wire this_vga_signals_M_vcounter_q_7;
    wire \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ;
    wire this_vga_signals_M_vcounter_q_8;
    wire \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ;
    wire \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ;
    wire \this_vga_signals.N_933_0 ;
    wire \this_vga_signals.N_1188_g ;
    wire N_422_2_cascade_;
    wire N_458_i;
    wire \this_vga_signals.M_vcounter_q_6_repZ0Z1 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_8 ;
    wire \this_vga_signals.M_vcounter_qZ0Z_9 ;
    wire \this_vga_signals.M_vcounter_q_fastZ0Z_7 ;
    wire \this_vga_signals.mult1_un40_sum_ac0_3_1_1 ;
    wire \this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3 ;
    wire \this_start_data_delay.N_424 ;
    wire M_this_spr_ram_write_data_0;
    wire M_this_state_qZ0Z_11;
    wire \this_start_data_delay.N_245_0_cascade_ ;
    wire un20_i_a4_0_a2_0_a2_1;
    wire M_this_state_qZ0Z_13;
    wire un20_i_a4_0_a2_2;
    wire N_241_0;
    wire \this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_ ;
    wire \this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0 ;
    wire M_this_state_qZ0Z_12;
    wire \this_start_data_delay.N_245_0 ;
    wire M_this_state_qZ0Z_7;
    wire M_this_state_qZ0Z_8;
    wire port_address_in_2;
    wire port_address_in_6;
    wire this_vga_signals_M_this_state_d28_0_a2_0_1;
    wire N_1264_0;
    wire \this_start_data_delay.N_387 ;
    wire port_address_in_0;
    wire port_address_in_4;
    wire \this_start_data_delay.N_337_cascade_ ;
    wire \this_start_data_delay.N_386 ;
    wire M_this_state_qZ0Z_6;
    wire M_this_state_qZ0Z_5;
    wire \this_start_data_delay.N_239_0 ;
    wire M_this_state_qZ0Z_3;
    wire M_this_state_qZ0Z_2;
    wire M_this_state_qZ0Z_1;
    wire \this_start_data_delay.N_420_3 ;
    wire \this_start_data_delay.N_23_1_0 ;
    wire \this_start_data_delay.N_344_cascade_ ;
    wire N_465;
    wire \this_start_data_delay.N_246_0 ;
    wire \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0 ;
    wire M_last_q_RNIE8SF1;
    wire M_this_ext_address_qZ0Z_0;
    wire bfn_21_24_0_;
    wire M_this_ext_address_qZ0Z_1;
    wire un1_M_this_ext_address_q_cry_0;
    wire M_this_ext_address_qZ0Z_2;
    wire un1_M_this_ext_address_q_cry_1;
    wire M_this_ext_address_qZ0Z_3;
    wire un1_M_this_ext_address_q_cry_2;
    wire M_this_ext_address_qZ0Z_4;
    wire un1_M_this_ext_address_q_cry_3;
    wire M_this_ext_address_qZ0Z_5;
    wire un1_M_this_ext_address_q_cry_4;
    wire M_this_ext_address_qZ0Z_6;
    wire un1_M_this_ext_address_q_cry_5;
    wire M_this_ext_address_qZ0Z_7;
    wire un1_M_this_ext_address_q_cry_6;
    wire un1_M_this_ext_address_q_cry_7;
    wire M_this_ext_address_qZ0Z_8;
    wire bfn_21_25_0_;
    wire M_this_ext_address_qZ0Z_9;
    wire un1_M_this_ext_address_q_cry_8;
    wire M_this_ext_address_qZ0Z_10;
    wire un1_M_this_ext_address_q_cry_9;
    wire M_this_ext_address_qZ0Z_11;
    wire un1_M_this_ext_address_q_cry_10;
    wire M_this_ext_address_qZ0Z_12;
    wire un1_M_this_ext_address_q_cry_11;
    wire M_this_ext_address_qZ0Z_13;
    wire un1_M_this_ext_address_q_cry_12;
    wire M_this_ext_address_qZ0Z_14;
    wire un1_M_this_ext_address_q_cry_13;
    wire N_295;
    wire un1_M_this_ext_address_q_cry_14;
    wire M_this_ext_address_qZ0Z_15;
    wire \this_start_data_delay.N_231_0 ;
    wire M_this_reset_cond_out_g_0;
    wire \this_start_data_delay.N_227_0 ;
    wire \this_start_data_delay.N_242_0 ;
    wire \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_ ;
    wire N_220_0;
    wire M_this_state_qZ0Z_10;
    wire N_930;
    wire M_this_state_qZ0Z_9;
    wire M_this_state_qZ0Z_4;
    wire \this_start_data_delay.N_332 ;
    wire port_data_c_0;
    wire M_this_map_ram_write_data_0;
    wire led_c_1;
    wire N_466;
    wire led_c_7;
    wire port_data_c_3;
    wire M_this_map_ram_write_data_3;
    wire port_data_c_1;
    wire M_this_map_ram_write_data_1;
    wire port_data_c_2;
    wire M_this_map_ram_write_data_2;
    wire port_data_c_4;
    wire M_this_map_ram_write_data_4;
    wire port_data_c_6;
    wire M_this_map_ram_write_data_6;
    wire port_data_c_5;
    wire M_this_map_ram_write_data_5;
    wire port_data_c_7;
    wire M_this_map_ram_write_data_7;
    wire M_this_state_d_0_sqmuxa;
    wire M_this_map_address_qZ0Z_0;
    wire bfn_26_25_0_;
    wire M_this_map_address_qZ0Z_1;
    wire un1_M_this_map_address_q_cry_0;
    wire M_this_map_address_qZ0Z_2;
    wire un1_M_this_map_address_q_cry_1;
    wire M_this_map_address_qZ0Z_3;
    wire un1_M_this_map_address_q_cry_2;
    wire M_this_map_address_qZ0Z_4;
    wire un1_M_this_map_address_q_cry_3;
    wire M_this_map_address_qZ0Z_5;
    wire un1_M_this_map_address_q_cry_4;
    wire M_this_map_address_qZ0Z_6;
    wire un1_M_this_map_address_q_cry_5;
    wire M_this_map_address_qZ0Z_7;
    wire un1_M_this_map_address_q_cry_6;
    wire un1_M_this_map_address_q_cry_7;
    wire M_this_map_address_qZ0Z_8;
    wire bfn_26_26_0_;
    wire N_93;
    wire un1_M_this_map_address_q_cry_8;
    wire M_this_map_address_qZ0Z_9;
    wire _gnd_net_;
    wire clk_0_c_g;
    wire N_527_g;

    defparam \this_map_ram.mem_mem_0_0_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_0_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,dangling_wire_1,M_this_map_ram_read_data_3,dangling_wire_2,dangling_wire_3,dangling_wire_4,M_this_map_ram_read_data_2,dangling_wire_5,dangling_wire_6,dangling_wire_7,M_this_map_ram_read_data_1,dangling_wire_8,dangling_wire_9,dangling_wire_10,M_this_map_ram_read_data_0,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__23300,N__22445,N__22505,N__22556,N__22613,N__25064,N__24110,N__24188,N__24266,N__24329}),
            .WADDR({dangling_wire_13,N__39461,N__39560,N__39590,N__39617,N__38375,N__38405,N__38432,N__38462,N__38492,N__38519}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__37772,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__37535,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__37658,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__38024,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__39418),
            .RE(N__25718),
            .WCLKE(N__38630),
            .WCLK(N__39419),
            .WE(N__25720));
    defparam \this_map_ram.mem_mem_0_1_physical .WRITE_MODE=2;
    defparam \this_map_ram.mem_mem_0_1_physical .READ_MODE=2;
    SB_RAM40_4K \this_map_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_42,dangling_wire_43,M_this_map_ram_read_data_7,dangling_wire_44,dangling_wire_45,dangling_wire_46,M_this_map_ram_read_data_6,dangling_wire_47,dangling_wire_48,dangling_wire_49,M_this_map_ram_read_data_5,dangling_wire_50,dangling_wire_51,dangling_wire_52,M_this_map_ram_read_data_4,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__23293,N__22439,N__22499,N__22546,N__22607,N__25058,N__24104,N__24182,N__24260,N__24319}),
            .WADDR({dangling_wire_55,N__39455,N__39554,N__39584,N__39611,N__38369,N__38399,N__38426,N__38456,N__38486,N__38513}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__38636,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__37259,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__38780,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__37406,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__39428),
            .RE(N__25719),
            .WCLKE(N__38625),
            .WCLK(N__39429),
            .WE(N__25721));
    defparam \this_oam_ram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_0_physical  (
            .RDATA({M_this_oam_ram_read_data_15,M_this_oam_ram_read_data_14,M_this_oam_ram_read_data_13,M_this_oam_ram_read_data_12,M_this_oam_ram_read_data_11,M_this_oam_ram_read_data_10,M_this_oam_ram_read_data_9,M_this_oam_ram_read_data_8,M_this_oam_ram_read_data_7,M_this_oam_ram_read_data_6,M_this_oam_ram_read_data_5,M_this_oam_ram_read_data_4,M_this_oam_ram_read_data_3,M_this_oam_ram_read_data_2,M_this_oam_ram_read_data_1,M_this_oam_ram_read_data_0}),
            .RADDR({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,N__18947,N__18680,N__18260,N__18349,N__18425,N__18551}),
            .WADDR({dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,N__17198,N__17231,N__19520,N__19481,N__19604,N__19568}),
            .MASK({dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .WDATA({N__15080,N__14846,N__15086,N__16637,N__17549,N__16649,N__17576,N__15038,N__15206,N__14978,N__15212,N__17567,N__15023,N__17594,N__17627,N__19229}),
            .RCLKE(),
            .RCLK(N__39431),
            .RE(N__25678),
            .WCLKE(N__19391),
            .WCLK(N__39432),
            .WE(N__25680));
    defparam \this_oam_ram.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_oam_ram.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_oam_ram.mem_mem_0_1_physical  (
            .RDATA({M_this_oam_ram_read_data_31,M_this_oam_ram_read_data_30,M_this_oam_ram_read_data_29,M_this_oam_ram_read_data_28,M_this_oam_ram_read_data_27,M_this_oam_ram_read_data_26,M_this_oam_ram_read_data_25,M_this_oam_ram_read_data_24,M_this_oam_ram_read_data_23,M_this_oam_ram_read_data_22,M_this_oam_ram_read_data_21,M_this_oam_ram_read_data_20,M_this_oam_ram_read_data_19,M_this_oam_ram_read_data_18,M_this_oam_ram_read_data_17,M_this_oam_ram_read_data_16}),
            .RADDR({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,N__18941,N__18674,N__18254,N__18336,N__18419,N__18545}),
            .WADDR({dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,N__17192,N__17225,N__19514,N__19475,N__19598,N__19562}),
            .MASK({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .WDATA({N__16601,N__15464,N__15452,N__17756,N__15470,N__19406,N__17747,N__15446,N__16790,N__15149,N__16802,N__17606,N__17768,N__15074,N__15458,N__15158}),
            .RCLKE(),
            .RCLK(N__39433),
            .RE(N__25679),
            .WCLKE(N__19390),
            .WCLK(N__39434),
            .WE(N__25681));
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_0_physical  (
            .RDATA({\this_ppu.oam_cache.mem_15 ,\this_ppu.oam_cache.mem_14 ,\this_ppu.oam_cache.mem_13 ,\this_ppu.oam_cache.mem_12 ,\this_ppu.oam_cache.mem_11 ,\this_ppu.oam_cache.mem_10 ,\this_ppu.oam_cache.mem_9 ,\this_ppu.oam_cache.mem_8 ,\this_ppu.oam_cache.mem_7 ,\this_ppu.oam_cache.mem_6 ,\this_ppu.oam_cache.mem_5 ,\this_ppu.oam_cache.mem_4 ,\this_ppu.oam_cache.mem_3 ,\this_ppu.oam_cache.mem_2 ,\this_ppu.oam_cache.mem_1 ,\this_ppu.oam_cache.mem_0 }),
            .RADDR({dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,N__18185,N__14735,N__14720,N__14699}),
            .WADDR({dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,N__13709,N__13412,N__13367,N__13454}),
            .MASK({dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165}),
            .WDATA({N__13295,N__13319,N__23783,N__23009,N__19181,N__13220,N__13238,N__13259,N__13631,N__13283,N__13655,N__13643,N__13289,N__13667,N__13619,N__13673}),
            .RCLKE(),
            .RCLK(N__39387),
            .RE(N__25503),
            .WCLKE(N__23950),
            .WCLK(N__39388),
            .WE(N__25599));
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \this_ppu.oam_cache.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,\this_ppu.oam_cache.mem_18 ,\this_ppu.oam_cache.mem_17 ,\this_ppu.oam_cache.mem_16 }),
            .RADDR({dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,N__18179,N__14729,N__14714,N__14693}),
            .WADDR({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,N__13701,N__13404,N__13361,N__13446}),
            .MASK({dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208}),
            .WDATA({N__15053,N__14831,N__15170,N__15191,N__23336,N__14855,N__14876,N__14903,N__14927,N__14750,N__14756,N__15101,N__15140,N__23369,N__23417,N__23459}),
            .RCLKE(),
            .RCLK(N__39400),
            .RE(N__25543),
            .WCLKE(N__24005),
            .WCLK(N__39401),
            .WE(N__25581));
    defparam \this_spr_ram.mem_mem_0_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,\this_spr_ram.mem_out_bus0_1 ,dangling_wire_213,dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,\this_spr_ram.mem_out_bus0_0 ,dangling_wire_220,dangling_wire_221,dangling_wire_222}),
            .RADDR({N__20314,N__20580,N__22983,N__32561,N__26290,N__15846,N__16008,N__17429,N__24483,N__24797,N__20147}),
            .WADDR({N__28912,N__29101,N__29349,N__29570,N__27113,N__27334,N__27521,N__27806,N__28049,N__28207,N__28414}),
            .MASK({dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238}),
            .WDATA({dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,N__32373,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,N__35085,dangling_wire_250,dangling_wire_251,dangling_wire_252}),
            .RCLKE(),
            .RCLK(N__39298),
            .RE(N__25722),
            .WCLKE(N__16753),
            .WCLK(N__39299),
            .WE(N__25724));
    defparam \this_spr_ram.mem_mem_0_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_0_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_0_1_physical  (
            .RDATA({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,\this_spr_ram.mem_out_bus0_3 ,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,\this_spr_ram.mem_out_bus0_2 ,dangling_wire_264,dangling_wire_265,dangling_wire_266}),
            .RADDR({N__20315,N__20581,N__22921,N__32535,N__26219,N__15827,N__16065,N__17455,N__24506,N__24738,N__20148}),
            .WADDR({N__28903,N__29100,N__29348,N__29569,N__27073,N__27280,N__27550,N__27802,N__28055,N__28236,N__28477}),
            .MASK({dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282}),
            .WDATA({dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__32818,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,N__34276,dangling_wire_294,dangling_wire_295,dangling_wire_296}),
            .RCLKE(),
            .RCLK(N__39291),
            .RE(N__25723),
            .WCLKE(N__16757),
            .WCLK(N__39292),
            .WE(N__25766));
    defparam \this_spr_ram.mem_mem_1_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_0_physical  (
            .RDATA({dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,\this_spr_ram.mem_out_bus1_1 ,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307,\this_spr_ram.mem_out_bus1_0 ,dangling_wire_308,dangling_wire_309,dangling_wire_310}),
            .RADDR({N__20350,N__20619,N__22993,N__32562,N__26289,N__15872,N__16088,N__17475,N__24501,N__24814,N__20176}),
            .WADDR({N__28902,N__29121,N__29354,N__29576,N__27130,N__27281,N__27497,N__27795,N__28048,N__28257,N__28495}),
            .MASK({dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326}),
            .WDATA({dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,N__32374,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__35097,dangling_wire_338,dangling_wire_339,dangling_wire_340}),
            .RCLKE(),
            .RCLK(N__39284),
            .RE(N__25795),
            .WCLKE(N__16774),
            .WCLK(N__39285),
            .WE(N__25580));
    defparam \this_spr_ram.mem_mem_1_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_1_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_1_1_physical  (
            .RDATA({dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,\this_spr_ram.mem_out_bus1_3 ,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,dangling_wire_351,\this_spr_ram.mem_out_bus1_2 ,dangling_wire_352,dangling_wire_353,dangling_wire_354}),
            .RADDR({N__20351,N__20620,N__22987,N__32563,N__26294,N__15873,N__16089,N__17489,N__24525,N__24801,N__20177}),
            .WADDR({N__28877,N__29028,N__29353,N__29575,N__27137,N__27282,N__27525,N__27775,N__28006,N__28269,N__28506}),
            .MASK({dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370}),
            .WDATA({dangling_wire_371,dangling_wire_372,dangling_wire_373,dangling_wire_374,N__32819,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,N__34282,dangling_wire_382,dangling_wire_383,dangling_wire_384}),
            .RCLKE(),
            .RCLK(N__39280),
            .RE(N__25796),
            .WCLKE(N__16778),
            .WCLK(N__39281),
            .WE(N__25797));
    defparam \this_spr_ram.mem_mem_2_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_0_physical  (
            .RDATA({dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,\this_spr_ram.mem_out_bus2_1 ,dangling_wire_389,dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,\this_spr_ram.mem_out_bus2_0 ,dangling_wire_396,dangling_wire_397,dangling_wire_398}),
            .RADDR({N__20405,N__20648,N__22994,N__32588,N__26263,N__15888,N__16109,N__17501,N__24536,N__24836,N__20146}),
            .WADDR({N__28868,N__29047,N__29286,N__29571,N__27134,N__27316,N__27566,N__27742,N__28005,N__28274,N__28505}),
            .MASK({dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414}),
            .WDATA({dangling_wire_415,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__32396,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,N__35102,dangling_wire_426,dangling_wire_427,dangling_wire_428}),
            .RCLKE(),
            .RCLK(N__39282),
            .RE(N__25800),
            .WCLKE(N__30722),
            .WCLK(N__39283),
            .WE(N__25799));
    defparam \this_spr_ram.mem_mem_2_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_2_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_2_1_physical  (
            .RDATA({dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,\this_spr_ram.mem_out_bus2_3 ,dangling_wire_433,dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,\this_spr_ram.mem_out_bus2_2 ,dangling_wire_440,dangling_wire_441,dangling_wire_442}),
            .RADDR({N__20401,N__20647,N__22989,N__32587,N__26300,N__15887,N__16108,N__17497,N__24502,N__24832,N__20145}),
            .WADDR({N__28869,N__29080,N__29341,N__29546,N__27120,N__27317,N__27496,N__27744,N__28050,N__28270,N__28491}),
            .MASK({dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458}),
            .WDATA({dangling_wire_459,dangling_wire_460,dangling_wire_461,dangling_wire_462,N__32814,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,N__34277,dangling_wire_470,dangling_wire_471,dangling_wire_472}),
            .RCLKE(),
            .RCLK(N__39286),
            .RE(N__25801),
            .WCLKE(N__30718),
            .WCLK(N__39287),
            .WE(N__25798));
    defparam \this_spr_ram.mem_mem_3_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_0_physical  (
            .RDATA({dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,\this_spr_ram.mem_out_bus3_1 ,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,\this_spr_ram.mem_out_bus3_0 ,dangling_wire_484,dangling_wire_485,dangling_wire_486}),
            .RADDR({N__20393,N__20640,N__22988,N__32580,N__26220,N__15856,N__16101,N__17490,N__24548,N__24739,N__20198}),
            .WADDR({N__28870,N__29081,N__29340,N__29550,N__27066,N__27319,N__27562,N__27743,N__28051,N__28262,N__28470}),
            .MASK({dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491,dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502}),
            .WDATA({dangling_wire_503,dangling_wire_504,dangling_wire_505,dangling_wire_506,N__32392,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,N__35098,dangling_wire_514,dangling_wire_515,dangling_wire_516}),
            .RCLKE(),
            .RCLK(N__39294),
            .RE(N__25777),
            .WCLKE(N__30113),
            .WCLK(N__39295),
            .WE(N__25788));
    defparam \this_spr_ram.mem_mem_3_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_3_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_3_1_physical  (
            .RDATA({dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,\this_spr_ram.mem_out_bus3_3 ,dangling_wire_521,dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,dangling_wire_526,dangling_wire_527,\this_spr_ram.mem_out_bus3_2 ,dangling_wire_528,dangling_wire_529,dangling_wire_530}),
            .RADDR({N__20379,N__20627,N__22972,N__32579,N__26295,N__15854,N__16046,N__17479,N__24544,N__24825,N__20192}),
            .WADDR({N__28900,N__29105,N__29311,N__29514,N__27106,N__27318,N__27555,N__27784,N__28031,N__28247,N__28469}),
            .MASK({dangling_wire_531,dangling_wire_532,dangling_wire_533,dangling_wire_534,dangling_wire_535,dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546}),
            .WDATA({dangling_wire_547,dangling_wire_548,dangling_wire_549,dangling_wire_550,N__32801,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,N__34263,dangling_wire_558,dangling_wire_559,dangling_wire_560}),
            .RCLKE(),
            .RCLK(N__39303),
            .RE(N__25776),
            .WCLKE(N__30109),
            .WCLK(N__39304),
            .WE(N__25787));
    defparam \this_spr_ram.mem_mem_4_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_0_physical  (
            .RDATA({dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,\this_spr_ram.mem_out_bus4_1 ,dangling_wire_565,dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,dangling_wire_570,dangling_wire_571,\this_spr_ram.mem_out_bus4_0 ,dangling_wire_572,dangling_wire_573,dangling_wire_574}),
            .RADDR({N__20359,N__20622,N__22971,N__32565,N__26296,N__15853,N__16091,N__17428,N__24537,N__24815,N__20178}),
            .WADDR({N__28901,N__29122,N__29318,N__29515,N__27079,N__27343,N__27540,N__27785,N__28004,N__28223,N__28437}),
            .MASK({dangling_wire_575,dangling_wire_576,dangling_wire_577,dangling_wire_578,dangling_wire_579,dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590}),
            .WDATA({dangling_wire_591,dangling_wire_592,dangling_wire_593,dangling_wire_594,N__32385,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,N__35089,dangling_wire_602,dangling_wire_603,dangling_wire_604}),
            .RCLKE(),
            .RCLK(N__39315),
            .RE(N__25737),
            .WCLKE(N__32246),
            .WCLK(N__39314),
            .WE(N__25765));
    defparam \this_spr_ram.mem_mem_4_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_4_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_4_1_physical  (
            .RDATA({dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,\this_spr_ram.mem_out_bus4_3 ,dangling_wire_609,dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,dangling_wire_614,dangling_wire_615,\this_spr_ram.mem_out_bus4_2 ,dangling_wire_616,dangling_wire_617,dangling_wire_618}),
            .RADDR({N__20322,N__20588,N__22941,N__32564,N__26276,N__15893,N__16090,N__17463,N__24526,N__24802,N__20119}),
            .WADDR({N__28911,N__29135,N__29285,N__29448,N__27033,N__27344,N__27463,N__27770,N__28037,N__28125,N__28429}),
            .MASK({dangling_wire_619,dangling_wire_620,dangling_wire_621,dangling_wire_622,dangling_wire_623,dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634}),
            .WDATA({dangling_wire_635,dangling_wire_636,dangling_wire_637,dangling_wire_638,N__32815,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,N__34245,dangling_wire_646,dangling_wire_647,dangling_wire_648}),
            .RCLKE(),
            .RCLK(N__39328),
            .RE(N__25736),
            .WCLKE(N__32245),
            .WCLK(N__39329),
            .WE(N__25764));
    defparam \this_spr_ram.mem_mem_5_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_0_physical  (
            .RDATA({dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,\this_spr_ram.mem_out_bus5_1 ,dangling_wire_653,dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,dangling_wire_658,dangling_wire_659,\this_spr_ram.mem_out_bus5_0 ,dangling_wire_660,dangling_wire_661,dangling_wire_662}),
            .RADDR({N__20352,N__20621,N__22940,N__32537,N__26279,N__15889,N__16073,N__17462,N__24510,N__24784,N__20155}),
            .WADDR({N__28898,N__29142,N__29287,N__29572,N__27074,N__27336,N__27533,N__27771,N__28036,N__28191,N__28430}),
            .MASK({dangling_wire_663,dangling_wire_664,dangling_wire_665,dangling_wire_666,dangling_wire_667,dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678}),
            .WDATA({dangling_wire_679,dangling_wire_680,dangling_wire_681,dangling_wire_682,N__32375,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,N__35072,dangling_wire_690,dangling_wire_691,dangling_wire_692}),
            .RCLKE(),
            .RCLK(N__39347),
            .RE(N__25683),
            .WCLKE(N__31837),
            .WCLK(N__39348),
            .WE(N__25684));
    defparam \this_spr_ram.mem_mem_5_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_5_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_5_1_physical  (
            .RDATA({dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,\this_spr_ram.mem_out_bus5_3 ,dangling_wire_697,dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,dangling_wire_702,dangling_wire_703,\this_spr_ram.mem_out_bus5_2 ,dangling_wire_704,dangling_wire_705,dangling_wire_706}),
            .RADDR({N__20377,N__20623,N__22900,N__32536,N__26277,N__15880,N__16072,N__17443,N__24462,N__24758,N__20165}),
            .WADDR({N__28899,N__29143,N__29288,N__29555,N__27075,N__27335,N__27553,N__27763,N__28032,N__28203,N__28465}),
            .MASK({dangling_wire_707,dangling_wire_708,dangling_wire_709,dangling_wire_710,dangling_wire_711,dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722}),
            .WDATA({dangling_wire_723,dangling_wire_724,dangling_wire_725,dangling_wire_726,N__32775,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,N__34244,dangling_wire_734,dangling_wire_735,dangling_wire_736}),
            .RCLKE(),
            .RCLK(N__39364),
            .RE(N__25685),
            .WCLKE(N__31838),
            .WCLK(N__39365),
            .WE(N__25717));
    defparam \this_spr_ram.mem_mem_6_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_0_physical  (
            .RDATA({dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,\this_spr_ram.mem_out_bus6_1 ,dangling_wire_741,dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,dangling_wire_746,dangling_wire_747,\this_spr_ram.mem_out_bus6_0 ,dangling_wire_748,dangling_wire_749,dangling_wire_750}),
            .RADDR({N__20378,N__20639,N__22859,N__32555,N__26278,N__15837,N__16047,N__17439,N__24443,N__24694,N__20185}),
            .WADDR({N__28894,N__29147,N__29289,N__29551,N__27105,N__27320,N__27554,N__27762,N__28052,N__28235,N__28490}),
            .MASK({dangling_wire_751,dangling_wire_752,dangling_wire_753,dangling_wire_754,dangling_wire_755,dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766}),
            .WDATA({dangling_wire_767,dangling_wire_768,dangling_wire_769,dangling_wire_770,N__32360,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,N__35051,dangling_wire_778,dangling_wire_779,dangling_wire_780}),
            .RCLKE(),
            .RCLK(N__39379),
            .RE(N__25618),
            .WCLKE(N__23557),
            .WCLK(N__39380),
            .WE(N__25625));
    defparam \this_spr_ram.mem_mem_6_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_6_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_6_1_physical  (
            .RDATA({dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,\this_spr_ram.mem_out_bus6_3 ,dangling_wire_785,dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,dangling_wire_790,dangling_wire_791,\this_spr_ram.mem_out_bus6_2 ,dangling_wire_792,dangling_wire_793,dangling_wire_794}),
            .RADDR({N__20343,N__20612,N__22957,N__32556,N__26298,N__15822,N__15975,N__17350,N__24480,N__24770,N__20169}),
            .WADDR({N__28890,N__29099,N__29350,N__29562,N__27083,N__27276,N__27551,N__27774,N__28041,N__28184,N__28459}),
            .MASK({dangling_wire_795,dangling_wire_796,dangling_wire_797,dangling_wire_798,dangling_wire_799,dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810}),
            .WDATA({dangling_wire_811,dangling_wire_812,dangling_wire_813,dangling_wire_814,N__32816,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,N__34278,dangling_wire_822,dangling_wire_823,dangling_wire_824}),
            .RCLKE(),
            .RCLK(N__39406),
            .RE(N__25544),
            .WCLKE(N__23564),
            .WCLK(N__39407),
            .WE(N__25582));
    defparam \this_spr_ram.mem_mem_7_0_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_0_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_0_physical  (
            .RDATA({dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,\this_spr_ram.mem_out_bus7_1 ,dangling_wire_829,dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,dangling_wire_834,dangling_wire_835,\this_spr_ram.mem_out_bus7_0 ,dangling_wire_836,dangling_wire_837,dangling_wire_838}),
            .RADDR({N__20389,N__20637,N__22967,N__32557,N__26299,N__15826,N__16006,N__17351,N__24481,N__24780,N__20196}),
            .WADDR({N__28913,N__29098,N__29351,N__29573,N__27135,N__27333,N__27552,N__27772,N__28054,N__28243,N__28507}),
            .MASK({dangling_wire_839,dangling_wire_840,dangling_wire_841,dangling_wire_842,dangling_wire_843,dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854}),
            .WDATA({dangling_wire_855,dangling_wire_856,dangling_wire_857,dangling_wire_858,N__32372,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,N__35096,dangling_wire_866,dangling_wire_867,dangling_wire_868}),
            .RCLKE(),
            .RCLK(N__39415),
            .RE(N__25660),
            .WCLKE(N__16714),
            .WCLK(N__39416),
            .WE(N__25601));
    defparam \this_spr_ram.mem_mem_7_1_physical .WRITE_MODE=3;
    defparam \this_spr_ram.mem_mem_7_1_physical .READ_MODE=3;
    SB_RAM40_4K \this_spr_ram.mem_mem_7_1_physical  (
            .RDATA({dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,\this_spr_ram.mem_out_bus7_3 ,dangling_wire_873,dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,dangling_wire_878,dangling_wire_879,\this_spr_ram.mem_out_bus7_2 ,dangling_wire_880,dangling_wire_881,dangling_wire_882}),
            .RADDR({N__20400,N__20638,N__22982,N__32578,N__26297,N__15855,N__16007,N__17374,N__24482,N__24796,N__20197}),
            .WADDR({N__28907,N__29120,N__29352,N__29574,N__27136,N__27312,N__27532,N__27773,N__28053,N__28261,N__28508}),
            .MASK({dangling_wire_883,dangling_wire_884,dangling_wire_885,dangling_wire_886,dangling_wire_887,dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898}),
            .WDATA({dangling_wire_899,dangling_wire_900,dangling_wire_901,dangling_wire_902,N__32817,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,N__34283,dangling_wire_910,dangling_wire_911,dangling_wire_912}),
            .RCLKE(),
            .RCLK(N__39425),
            .RE(N__25661),
            .WCLKE(N__16721),
            .WCLK(N__39426),
            .WE(N__25602));
    defparam \this_vram.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \this_vram.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \this_vram.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917,dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,dangling_wire_922,dangling_wire_923,dangling_wire_924,M_this_vram_read_data_3,M_this_vram_read_data_2,M_this_vram_read_data_1,M_this_vram_read_data_0}),
            .RADDR({dangling_wire_925,dangling_wire_926,dangling_wire_927,N__26426,N__12728,N__13154,N__13127,N__13169,N__13019,N__12839,N__12983}),
            .WADDR({dangling_wire_928,dangling_wire_929,dangling_wire_930,N__23264,N__17003,N__17027,N__16844,N__17897,N__16904,N__16976,N__16946}),
            .MASK({dangling_wire_931,dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,dangling_wire_943,dangling_wire_944,dangling_wire_945,dangling_wire_946}),
            .WDATA({dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,N__17786,N__18692,N__17846,N__16694}),
            .RCLKE(),
            .RCLK(N__39372),
            .RE(N__25515),
            .WCLKE(N__20930),
            .WCLK(N__39373),
            .WE(N__25600));
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__40095),
            .GLOBALBUFFEROUTPUT(clk_0_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__40097),
            .DIN(N__40096),
            .DOUT(N__40095),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__40097),
            .PADOUT(N__40096),
            .PADIN(N__40095),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_0_iopad (
            .OE(N__40086),
            .DIN(N__40085),
            .DOUT(N__40084),
            .PACKAGEPIN(debug[0]));
    defparam debug_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_0_preio (
            .PADOEN(N__40086),
            .PADOUT(N__40085),
            .PADIN(N__40084),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD debug_obuf_1_iopad (
            .OE(N__40077),
            .DIN(N__40076),
            .DOUT(N__40075),
            .PACKAGEPIN(debug[1]));
    defparam debug_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam debug_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO debug_obuf_1_preio (
            .PADOEN(N__40077),
            .PADOUT(N__40076),
            .PADIN(N__40075),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hblank_obuf_iopad (
            .OE(N__40068),
            .DIN(N__40067),
            .DOUT(N__40066),
            .PACKAGEPIN(hblank));
    defparam hblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hblank_obuf_preio (
            .PADOEN(N__40068),
            .PADOUT(N__40067),
            .PADIN(N__40066),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12920),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD hsync_obuf_iopad (
            .OE(N__40059),
            .DIN(N__40058),
            .DOUT(N__40057),
            .PACKAGEPIN(hsync));
    defparam hsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam hsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO hsync_obuf_preio (
            .PADOEN(N__40059),
            .PADOUT(N__40058),
            .PADIN(N__40057),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12935),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_0_iopad (
            .OE(N__40050),
            .DIN(N__40049),
            .DOUT(N__40048),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__40050),
            .PADOUT(N__40049),
            .PADIN(N__40048),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__25805),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_1_iopad (
            .OE(N__40041),
            .DIN(N__40040),
            .DOUT(N__40039),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__40041),
            .PADOUT(N__40040),
            .PADIN(N__40039),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__38012),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_2_iopad (
            .OE(N__40032),
            .DIN(N__40031),
            .DOUT(N__40030),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__40032),
            .PADOUT(N__40031),
            .PADIN(N__40030),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_3_iopad (
            .OE(N__40023),
            .DIN(N__40022),
            .DOUT(N__40021),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__40023),
            .PADOUT(N__40022),
            .PADIN(N__40021),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_4_iopad (
            .OE(N__40014),
            .DIN(N__40013),
            .DOUT(N__40012),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__40014),
            .PADOUT(N__40013),
            .PADIN(N__40012),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_5_iopad (
            .OE(N__40005),
            .DIN(N__40004),
            .DOUT(N__40003),
            .PACKAGEPIN(led[5]));
    defparam led_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_5_preio (
            .PADOEN(N__40005),
            .PADOUT(N__40004),
            .PADIN(N__40003),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_6_iopad (
            .OE(N__39996),
            .DIN(N__39995),
            .DOUT(N__39994),
            .PACKAGEPIN(led[6]));
    defparam led_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_6_preio (
            .PADOEN(N__39996),
            .PADOUT(N__39995),
            .PADIN(N__39994),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34400),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD led_obuf_7_iopad (
            .OE(N__39987),
            .DIN(N__39986),
            .DOUT(N__39985),
            .PACKAGEPIN(led[7]));
    defparam led_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_7_preio (
            .PADOEN(N__39987),
            .PADOUT(N__39986),
            .PADIN(N__39985),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37913),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_address_iobuf_0_iopad (
            .OE(N__39978),
            .DIN(N__39977),
            .DOUT(N__39976),
            .PACKAGEPIN(port_address[0]));
    defparam port_address_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_0_preio (
            .PADOEN(N__39978),
            .PADOUT(N__39977),
            .PADIN(N__39976),
            .CLOCKENABLE(),
            .DIN0(port_address_in_0),
            .DIN1(),
            .DOUT0(N__35858),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15372));
    IO_PAD port_address_iobuf_1_iopad (
            .OE(N__39969),
            .DIN(N__39968),
            .DOUT(N__39967),
            .PACKAGEPIN(port_address[1]));
    defparam port_address_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_1_preio (
            .PADOEN(N__39969),
            .PADOUT(N__39968),
            .PADIN(N__39967),
            .CLOCKENABLE(),
            .DIN0(port_address_in_1),
            .DIN1(),
            .DOUT0(N__35840),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15404));
    IO_PAD port_address_iobuf_2_iopad (
            .OE(N__39960),
            .DIN(N__39959),
            .DOUT(N__39958),
            .PACKAGEPIN(port_address[2]));
    defparam port_address_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_2_preio (
            .PADOEN(N__39960),
            .PADOUT(N__39959),
            .PADIN(N__39958),
            .CLOCKENABLE(),
            .DIN0(port_address_in_2),
            .DIN1(),
            .DOUT0(N__36392),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15362));
    IO_PAD port_address_iobuf_3_iopad (
            .OE(N__39951),
            .DIN(N__39950),
            .DOUT(N__39949),
            .PACKAGEPIN(port_address[3]));
    defparam port_address_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_3_preio (
            .PADOEN(N__39951),
            .PADOUT(N__39950),
            .PADIN(N__39949),
            .CLOCKENABLE(),
            .DIN0(port_address_in_3),
            .DIN1(),
            .DOUT0(N__36368),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15440));
    IO_PAD port_address_iobuf_4_iopad (
            .OE(N__39942),
            .DIN(N__39941),
            .DOUT(N__39940),
            .PACKAGEPIN(port_address[4]));
    defparam port_address_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_4_preio (
            .PADOEN(N__39942),
            .PADOUT(N__39941),
            .PADIN(N__39940),
            .CLOCKENABLE(),
            .DIN0(port_address_in_4),
            .DIN1(),
            .DOUT0(N__36341),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15435));
    IO_PAD port_address_iobuf_5_iopad (
            .OE(N__39933),
            .DIN(N__39932),
            .DOUT(N__39931),
            .PACKAGEPIN(port_address[5]));
    defparam port_address_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_5_preio (
            .PADOEN(N__39933),
            .PADOUT(N__39932),
            .PADIN(N__39931),
            .CLOCKENABLE(),
            .DIN0(port_address_in_5),
            .DIN1(),
            .DOUT0(N__36314),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15424));
    IO_PAD port_address_iobuf_6_iopad (
            .OE(N__39924),
            .DIN(N__39923),
            .DOUT(N__39922),
            .PACKAGEPIN(port_address[6]));
    defparam port_address_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_6_preio (
            .PADOEN(N__39924),
            .PADOUT(N__39923),
            .PADIN(N__39922),
            .CLOCKENABLE(),
            .DIN0(port_address_in_6),
            .DIN1(),
            .DOUT0(N__36287),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15409));
    IO_PAD port_address_iobuf_7_iopad (
            .OE(N__39915),
            .DIN(N__39914),
            .DOUT(N__39913),
            .PACKAGEPIN(port_address[7]));
    defparam port_address_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_address_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_iobuf_7_preio (
            .PADOEN(N__39915),
            .PADOUT(N__39914),
            .PADIN(N__39913),
            .CLOCKENABLE(),
            .DIN0(port_address_in_7),
            .DIN1(),
            .DOUT0(N__36257),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15373));
    IO_PAD port_address_obuft_10_iopad (
            .OE(N__39906),
            .DIN(N__39905),
            .DOUT(N__39904),
            .PACKAGEPIN(port_address[10]));
    defparam port_address_obuft_10_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_10_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_10_preio (
            .PADOEN(N__39906),
            .PADOUT(N__39905),
            .PADIN(N__39904),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37250),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15364));
    IO_PAD port_address_obuft_11_iopad (
            .OE(N__39897),
            .DIN(N__39896),
            .DOUT(N__39895),
            .PACKAGEPIN(port_address[11]));
    defparam port_address_obuft_11_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_11_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_11_preio (
            .PADOEN(N__39897),
            .PADOUT(N__39896),
            .PADIN(N__39895),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37223),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15423));
    IO_PAD port_address_obuft_12_iopad (
            .OE(N__39888),
            .DIN(N__39887),
            .DOUT(N__39886),
            .PACKAGEPIN(port_address[12]));
    defparam port_address_obuft_12_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_12_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_12_preio (
            .PADOEN(N__39888),
            .PADOUT(N__39887),
            .PADIN(N__39886),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37190),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15436));
    IO_PAD port_address_obuft_13_iopad (
            .OE(N__39879),
            .DIN(N__39878),
            .DOUT(N__39877),
            .PACKAGEPIN(port_address[13]));
    defparam port_address_obuft_13_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_13_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_13_preio (
            .PADOEN(N__39879),
            .PADOUT(N__39878),
            .PADIN(N__39877),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37160),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15425));
    IO_PAD port_address_obuft_14_iopad (
            .OE(N__39870),
            .DIN(N__39869),
            .DOUT(N__39868),
            .PACKAGEPIN(port_address[14]));
    defparam port_address_obuft_14_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_14_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_14_preio (
            .PADOEN(N__39870),
            .PADOUT(N__39869),
            .PADIN(N__39868),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37130),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15408));
    IO_PAD port_address_obuft_15_iopad (
            .OE(N__39861),
            .DIN(N__39860),
            .DOUT(N__39859),
            .PACKAGEPIN(port_address[15]));
    defparam port_address_obuft_15_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_15_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_15_preio (
            .PADOEN(N__39861),
            .PADOUT(N__39860),
            .PADIN(N__39859),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37019),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15311));
    IO_PAD port_address_obuft_8_iopad (
            .OE(N__39852),
            .DIN(N__39851),
            .DOUT(N__39850),
            .PACKAGEPIN(port_address[8]));
    defparam port_address_obuft_8_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_8_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_8_preio (
            .PADOEN(N__39852),
            .PADOUT(N__39851),
            .PADIN(N__39850),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36227),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15363));
    IO_PAD port_address_obuft_9_iopad (
            .OE(N__39843),
            .DIN(N__39842),
            .DOUT(N__39841),
            .PACKAGEPIN(port_address[9]));
    defparam port_address_obuft_9_preio.NEG_TRIGGER=1'b0;
    defparam port_address_obuft_9_preio.PIN_TYPE=6'b101001;
    PRE_IO port_address_obuft_9_preio (
            .PADOEN(N__39843),
            .PADOUT(N__39842),
            .PADIN(N__39841),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__36197),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15403));
    IO_PAD port_clk_ibuf_iopad (
            .OE(N__39834),
            .DIN(N__39833),
            .DOUT(N__39832),
            .PACKAGEPIN(port_clk));
    defparam port_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_clk_ibuf_preio (
            .PADOEN(N__39834),
            .PADOUT(N__39833),
            .PADIN(N__39832),
            .CLOCKENABLE(),
            .DIN0(port_clk_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_0_iopad (
            .OE(N__39825),
            .DIN(N__39824),
            .DOUT(N__39823),
            .PACKAGEPIN(port_data[0]));
    defparam port_data_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_0_preio (
            .PADOEN(N__39825),
            .PADOUT(N__39824),
            .PADIN(N__39823),
            .CLOCKENABLE(),
            .DIN0(port_data_c_0),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_1_iopad (
            .OE(N__39816),
            .DIN(N__39815),
            .DOUT(N__39814),
            .PACKAGEPIN(port_data[1]));
    defparam port_data_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_1_preio (
            .PADOEN(N__39816),
            .PADOUT(N__39815),
            .PADIN(N__39814),
            .CLOCKENABLE(),
            .DIN0(port_data_c_1),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_2_iopad (
            .OE(N__39807),
            .DIN(N__39806),
            .DOUT(N__39805),
            .PACKAGEPIN(port_data[2]));
    defparam port_data_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_2_preio (
            .PADOEN(N__39807),
            .PADOUT(N__39806),
            .PADIN(N__39805),
            .CLOCKENABLE(),
            .DIN0(port_data_c_2),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_3_iopad (
            .OE(N__39798),
            .DIN(N__39797),
            .DOUT(N__39796),
            .PACKAGEPIN(port_data[3]));
    defparam port_data_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_3_preio (
            .PADOEN(N__39798),
            .PADOUT(N__39797),
            .PADIN(N__39796),
            .CLOCKENABLE(),
            .DIN0(port_data_c_3),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_4_iopad (
            .OE(N__39789),
            .DIN(N__39788),
            .DOUT(N__39787),
            .PACKAGEPIN(port_data[4]));
    defparam port_data_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_4_preio (
            .PADOEN(N__39789),
            .PADOUT(N__39788),
            .PADIN(N__39787),
            .CLOCKENABLE(),
            .DIN0(port_data_c_4),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_5_iopad (
            .OE(N__39780),
            .DIN(N__39779),
            .DOUT(N__39778),
            .PACKAGEPIN(port_data[5]));
    defparam port_data_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_5_preio (
            .PADOEN(N__39780),
            .PADOUT(N__39779),
            .PADIN(N__39778),
            .CLOCKENABLE(),
            .DIN0(port_data_c_5),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_6_iopad (
            .OE(N__39771),
            .DIN(N__39770),
            .DOUT(N__39769),
            .PACKAGEPIN(port_data[6]));
    defparam port_data_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_6_preio (
            .PADOEN(N__39771),
            .PADOUT(N__39770),
            .PADIN(N__39769),
            .CLOCKENABLE(),
            .DIN0(port_data_c_6),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_ibuf_7_iopad (
            .OE(N__39762),
            .DIN(N__39761),
            .DOUT(N__39760),
            .PACKAGEPIN(port_data[7]));
    defparam port_data_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam port_data_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO port_data_ibuf_7_preio (
            .PADOEN(N__39762),
            .PADOUT(N__39761),
            .PADIN(N__39760),
            .CLOCKENABLE(),
            .DIN0(port_data_c_7),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_data_rw_obuf_iopad (
            .OE(N__39753),
            .DIN(N__39752),
            .DOUT(N__39751),
            .PACKAGEPIN(port_data_rw));
    defparam port_data_rw_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_data_rw_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_data_rw_obuf_preio (
            .PADOEN(N__39753),
            .PADOUT(N__39752),
            .PADIN(N__39751),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12716),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_dmab_obuf_iopad (
            .OE(N__39744),
            .DIN(N__39743),
            .DOUT(N__39742),
            .PACKAGEPIN(port_dmab));
    defparam port_dmab_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_dmab_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_dmab_obuf_preio (
            .PADOEN(N__39744),
            .PADOUT(N__39743),
            .PADIN(N__39742),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__34177),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_enb_ibuf_iopad (
            .OE(N__39735),
            .DIN(N__39734),
            .DOUT(N__39733),
            .PACKAGEPIN(port_enb));
    defparam port_enb_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam port_enb_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO port_enb_ibuf_preio (
            .PADOEN(N__39735),
            .PADOUT(N__39734),
            .PADIN(N__39733),
            .CLOCKENABLE(),
            .DIN0(port_enb_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_nmib_obuf_iopad (
            .OE(N__39726),
            .DIN(N__39725),
            .DOUT(N__39724),
            .PACKAGEPIN(port_nmib));
    defparam port_nmib_obuf_preio.NEG_TRIGGER=1'b0;
    defparam port_nmib_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO port_nmib_obuf_preio (
            .PADOEN(N__39726),
            .PADOUT(N__39725),
            .PADIN(N__39724),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__26387),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD port_rw_iobuf_iopad (
            .OE(N__39717),
            .DIN(N__39716),
            .DOUT(N__39715),
            .PACKAGEPIN(port_rw));
    defparam port_rw_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam port_rw_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO port_rw_iobuf_preio (
            .PADOEN(N__39717),
            .PADOUT(N__39716),
            .PADIN(N__39715),
            .CLOCKENABLE(),
            .DIN0(port_rw_in),
            .DIN1(),
            .DOUT0(N__25682),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__15352));
    IO_PAD rgb_obuf_0_iopad (
            .OE(N__39708),
            .DIN(N__39707),
            .DOUT(N__39706),
            .PACKAGEPIN(rgb[0]));
    defparam rgb_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_0_preio (
            .PADOEN(N__39708),
            .PADOUT(N__39707),
            .PADIN(N__39706),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12890),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_1_iopad (
            .OE(N__39699),
            .DIN(N__39698),
            .DOUT(N__39697),
            .PACKAGEPIN(rgb[1]));
    defparam rgb_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_1_preio (
            .PADOEN(N__39699),
            .PADOUT(N__39698),
            .PADIN(N__39697),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12791),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_2_iopad (
            .OE(N__39690),
            .DIN(N__39689),
            .DOUT(N__39688),
            .PACKAGEPIN(rgb[2]));
    defparam rgb_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_2_preio (
            .PADOEN(N__39690),
            .PADOUT(N__39689),
            .PADIN(N__39688),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12770),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_3_iopad (
            .OE(N__39681),
            .DIN(N__39680),
            .DOUT(N__39679),
            .PACKAGEPIN(rgb[3]));
    defparam rgb_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_3_preio (
            .PADOEN(N__39681),
            .PADOUT(N__39680),
            .PADIN(N__39679),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12809),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_4_iopad (
            .OE(N__39672),
            .DIN(N__39671),
            .DOUT(N__39670),
            .PACKAGEPIN(rgb[4]));
    defparam rgb_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_4_preio (
            .PADOEN(N__39672),
            .PADOUT(N__39671),
            .PADIN(N__39670),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12761),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rgb_obuf_5_iopad (
            .OE(N__39663),
            .DIN(N__39662),
            .DOUT(N__39661),
            .PACKAGEPIN(rgb[5]));
    defparam rgb_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam rgb_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO rgb_obuf_5_preio (
            .PADOEN(N__39663),
            .PADOUT(N__39662),
            .PADIN(N__39661),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12743),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__39654),
            .DIN(N__39653),
            .DOUT(N__39652),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__39654),
            .PADOUT(N__39653),
            .PADIN(N__39652),
            .CLOCKENABLE(),
            .DIN0(rst_n_c),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vblank_obuf_iopad (
            .OE(N__39645),
            .DIN(N__39644),
            .DOUT(N__39643),
            .PACKAGEPIN(vblank));
    defparam vblank_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vblank_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vblank_obuf_preio (
            .PADOEN(N__39645),
            .PADOUT(N__39644),
            .PADIN(N__39643),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__12899),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    IO_PAD vsync_obuf_iopad (
            .OE(N__39636),
            .DIN(N__39635),
            .DOUT(N__39634),
            .PACKAGEPIN(vsync));
    defparam vsync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam vsync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO vsync_obuf_preio (
            .PADOEN(N__39636),
            .PADOUT(N__39635),
            .PADIN(N__39634),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__29879),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    CascadeMux I__9910 (
            .O(N__39617),
            .I(N__39614));
    CascadeBuf I__9909 (
            .O(N__39614),
            .I(N__39611));
    CascadeMux I__9908 (
            .O(N__39611),
            .I(N__39608));
    InMux I__9907 (
            .O(N__39608),
            .I(N__39604));
    InMux I__9906 (
            .O(N__39607),
            .I(N__39601));
    LocalMux I__9905 (
            .O(N__39604),
            .I(N__39598));
    LocalMux I__9904 (
            .O(N__39601),
            .I(M_this_map_address_qZ0Z_6));
    Odrv4 I__9903 (
            .O(N__39598),
            .I(M_this_map_address_qZ0Z_6));
    InMux I__9902 (
            .O(N__39593),
            .I(un1_M_this_map_address_q_cry_5));
    CascadeMux I__9901 (
            .O(N__39590),
            .I(N__39587));
    CascadeBuf I__9900 (
            .O(N__39587),
            .I(N__39584));
    CascadeMux I__9899 (
            .O(N__39584),
            .I(N__39581));
    InMux I__9898 (
            .O(N__39581),
            .I(N__39578));
    LocalMux I__9897 (
            .O(N__39578),
            .I(N__39574));
    InMux I__9896 (
            .O(N__39577),
            .I(N__39571));
    Span4Mux_h I__9895 (
            .O(N__39574),
            .I(N__39568));
    LocalMux I__9894 (
            .O(N__39571),
            .I(M_this_map_address_qZ0Z_7));
    Odrv4 I__9893 (
            .O(N__39568),
            .I(M_this_map_address_qZ0Z_7));
    InMux I__9892 (
            .O(N__39563),
            .I(un1_M_this_map_address_q_cry_6));
    CascadeMux I__9891 (
            .O(N__39560),
            .I(N__39557));
    CascadeBuf I__9890 (
            .O(N__39557),
            .I(N__39554));
    CascadeMux I__9889 (
            .O(N__39554),
            .I(N__39551));
    InMux I__9888 (
            .O(N__39551),
            .I(N__39548));
    LocalMux I__9887 (
            .O(N__39548),
            .I(N__39544));
    InMux I__9886 (
            .O(N__39547),
            .I(N__39541));
    Span4Mux_h I__9885 (
            .O(N__39544),
            .I(N__39538));
    LocalMux I__9884 (
            .O(N__39541),
            .I(M_this_map_address_qZ0Z_8));
    Odrv4 I__9883 (
            .O(N__39538),
            .I(M_this_map_address_qZ0Z_8));
    InMux I__9882 (
            .O(N__39533),
            .I(bfn_26_26_0_));
    CascadeMux I__9881 (
            .O(N__39530),
            .I(N__39527));
    InMux I__9880 (
            .O(N__39527),
            .I(N__39514));
    InMux I__9879 (
            .O(N__39526),
            .I(N__39509));
    InMux I__9878 (
            .O(N__39525),
            .I(N__39509));
    InMux I__9877 (
            .O(N__39524),
            .I(N__39500));
    InMux I__9876 (
            .O(N__39523),
            .I(N__39500));
    InMux I__9875 (
            .O(N__39522),
            .I(N__39500));
    InMux I__9874 (
            .O(N__39521),
            .I(N__39500));
    InMux I__9873 (
            .O(N__39520),
            .I(N__39491));
    InMux I__9872 (
            .O(N__39519),
            .I(N__39491));
    InMux I__9871 (
            .O(N__39518),
            .I(N__39491));
    InMux I__9870 (
            .O(N__39517),
            .I(N__39491));
    LocalMux I__9869 (
            .O(N__39514),
            .I(N__39488));
    LocalMux I__9868 (
            .O(N__39509),
            .I(N__39481));
    LocalMux I__9867 (
            .O(N__39500),
            .I(N__39481));
    LocalMux I__9866 (
            .O(N__39491),
            .I(N__39481));
    Span4Mux_v I__9865 (
            .O(N__39488),
            .I(N__39478));
    Span4Mux_v I__9864 (
            .O(N__39481),
            .I(N__39475));
    Span4Mux_h I__9863 (
            .O(N__39478),
            .I(N__39472));
    Span4Mux_h I__9862 (
            .O(N__39475),
            .I(N__39469));
    Odrv4 I__9861 (
            .O(N__39472),
            .I(N_93));
    Odrv4 I__9860 (
            .O(N__39469),
            .I(N_93));
    InMux I__9859 (
            .O(N__39464),
            .I(un1_M_this_map_address_q_cry_8));
    CascadeMux I__9858 (
            .O(N__39461),
            .I(N__39458));
    CascadeBuf I__9857 (
            .O(N__39458),
            .I(N__39455));
    CascadeMux I__9856 (
            .O(N__39455),
            .I(N__39452));
    InMux I__9855 (
            .O(N__39452),
            .I(N__39449));
    LocalMux I__9854 (
            .O(N__39449),
            .I(N__39445));
    InMux I__9853 (
            .O(N__39448),
            .I(N__39442));
    Span4Mux_h I__9852 (
            .O(N__39445),
            .I(N__39439));
    LocalMux I__9851 (
            .O(N__39442),
            .I(M_this_map_address_qZ0Z_9));
    Odrv4 I__9850 (
            .O(N__39439),
            .I(M_this_map_address_qZ0Z_9));
    ClkMux I__9849 (
            .O(N__39434),
            .I(N__38969));
    ClkMux I__9848 (
            .O(N__39433),
            .I(N__38969));
    ClkMux I__9847 (
            .O(N__39432),
            .I(N__38969));
    ClkMux I__9846 (
            .O(N__39431),
            .I(N__38969));
    ClkMux I__9845 (
            .O(N__39430),
            .I(N__38969));
    ClkMux I__9844 (
            .O(N__39429),
            .I(N__38969));
    ClkMux I__9843 (
            .O(N__39428),
            .I(N__38969));
    ClkMux I__9842 (
            .O(N__39427),
            .I(N__38969));
    ClkMux I__9841 (
            .O(N__39426),
            .I(N__38969));
    ClkMux I__9840 (
            .O(N__39425),
            .I(N__38969));
    ClkMux I__9839 (
            .O(N__39424),
            .I(N__38969));
    ClkMux I__9838 (
            .O(N__39423),
            .I(N__38969));
    ClkMux I__9837 (
            .O(N__39422),
            .I(N__38969));
    ClkMux I__9836 (
            .O(N__39421),
            .I(N__38969));
    ClkMux I__9835 (
            .O(N__39420),
            .I(N__38969));
    ClkMux I__9834 (
            .O(N__39419),
            .I(N__38969));
    ClkMux I__9833 (
            .O(N__39418),
            .I(N__38969));
    ClkMux I__9832 (
            .O(N__39417),
            .I(N__38969));
    ClkMux I__9831 (
            .O(N__39416),
            .I(N__38969));
    ClkMux I__9830 (
            .O(N__39415),
            .I(N__38969));
    ClkMux I__9829 (
            .O(N__39414),
            .I(N__38969));
    ClkMux I__9828 (
            .O(N__39413),
            .I(N__38969));
    ClkMux I__9827 (
            .O(N__39412),
            .I(N__38969));
    ClkMux I__9826 (
            .O(N__39411),
            .I(N__38969));
    ClkMux I__9825 (
            .O(N__39410),
            .I(N__38969));
    ClkMux I__9824 (
            .O(N__39409),
            .I(N__38969));
    ClkMux I__9823 (
            .O(N__39408),
            .I(N__38969));
    ClkMux I__9822 (
            .O(N__39407),
            .I(N__38969));
    ClkMux I__9821 (
            .O(N__39406),
            .I(N__38969));
    ClkMux I__9820 (
            .O(N__39405),
            .I(N__38969));
    ClkMux I__9819 (
            .O(N__39404),
            .I(N__38969));
    ClkMux I__9818 (
            .O(N__39403),
            .I(N__38969));
    ClkMux I__9817 (
            .O(N__39402),
            .I(N__38969));
    ClkMux I__9816 (
            .O(N__39401),
            .I(N__38969));
    ClkMux I__9815 (
            .O(N__39400),
            .I(N__38969));
    ClkMux I__9814 (
            .O(N__39399),
            .I(N__38969));
    ClkMux I__9813 (
            .O(N__39398),
            .I(N__38969));
    ClkMux I__9812 (
            .O(N__39397),
            .I(N__38969));
    ClkMux I__9811 (
            .O(N__39396),
            .I(N__38969));
    ClkMux I__9810 (
            .O(N__39395),
            .I(N__38969));
    ClkMux I__9809 (
            .O(N__39394),
            .I(N__38969));
    ClkMux I__9808 (
            .O(N__39393),
            .I(N__38969));
    ClkMux I__9807 (
            .O(N__39392),
            .I(N__38969));
    ClkMux I__9806 (
            .O(N__39391),
            .I(N__38969));
    ClkMux I__9805 (
            .O(N__39390),
            .I(N__38969));
    ClkMux I__9804 (
            .O(N__39389),
            .I(N__38969));
    ClkMux I__9803 (
            .O(N__39388),
            .I(N__38969));
    ClkMux I__9802 (
            .O(N__39387),
            .I(N__38969));
    ClkMux I__9801 (
            .O(N__39386),
            .I(N__38969));
    ClkMux I__9800 (
            .O(N__39385),
            .I(N__38969));
    ClkMux I__9799 (
            .O(N__39384),
            .I(N__38969));
    ClkMux I__9798 (
            .O(N__39383),
            .I(N__38969));
    ClkMux I__9797 (
            .O(N__39382),
            .I(N__38969));
    ClkMux I__9796 (
            .O(N__39381),
            .I(N__38969));
    ClkMux I__9795 (
            .O(N__39380),
            .I(N__38969));
    ClkMux I__9794 (
            .O(N__39379),
            .I(N__38969));
    ClkMux I__9793 (
            .O(N__39378),
            .I(N__38969));
    ClkMux I__9792 (
            .O(N__39377),
            .I(N__38969));
    ClkMux I__9791 (
            .O(N__39376),
            .I(N__38969));
    ClkMux I__9790 (
            .O(N__39375),
            .I(N__38969));
    ClkMux I__9789 (
            .O(N__39374),
            .I(N__38969));
    ClkMux I__9788 (
            .O(N__39373),
            .I(N__38969));
    ClkMux I__9787 (
            .O(N__39372),
            .I(N__38969));
    ClkMux I__9786 (
            .O(N__39371),
            .I(N__38969));
    ClkMux I__9785 (
            .O(N__39370),
            .I(N__38969));
    ClkMux I__9784 (
            .O(N__39369),
            .I(N__38969));
    ClkMux I__9783 (
            .O(N__39368),
            .I(N__38969));
    ClkMux I__9782 (
            .O(N__39367),
            .I(N__38969));
    ClkMux I__9781 (
            .O(N__39366),
            .I(N__38969));
    ClkMux I__9780 (
            .O(N__39365),
            .I(N__38969));
    ClkMux I__9779 (
            .O(N__39364),
            .I(N__38969));
    ClkMux I__9778 (
            .O(N__39363),
            .I(N__38969));
    ClkMux I__9777 (
            .O(N__39362),
            .I(N__38969));
    ClkMux I__9776 (
            .O(N__39361),
            .I(N__38969));
    ClkMux I__9775 (
            .O(N__39360),
            .I(N__38969));
    ClkMux I__9774 (
            .O(N__39359),
            .I(N__38969));
    ClkMux I__9773 (
            .O(N__39358),
            .I(N__38969));
    ClkMux I__9772 (
            .O(N__39357),
            .I(N__38969));
    ClkMux I__9771 (
            .O(N__39356),
            .I(N__38969));
    ClkMux I__9770 (
            .O(N__39355),
            .I(N__38969));
    ClkMux I__9769 (
            .O(N__39354),
            .I(N__38969));
    ClkMux I__9768 (
            .O(N__39353),
            .I(N__38969));
    ClkMux I__9767 (
            .O(N__39352),
            .I(N__38969));
    ClkMux I__9766 (
            .O(N__39351),
            .I(N__38969));
    ClkMux I__9765 (
            .O(N__39350),
            .I(N__38969));
    ClkMux I__9764 (
            .O(N__39349),
            .I(N__38969));
    ClkMux I__9763 (
            .O(N__39348),
            .I(N__38969));
    ClkMux I__9762 (
            .O(N__39347),
            .I(N__38969));
    ClkMux I__9761 (
            .O(N__39346),
            .I(N__38969));
    ClkMux I__9760 (
            .O(N__39345),
            .I(N__38969));
    ClkMux I__9759 (
            .O(N__39344),
            .I(N__38969));
    ClkMux I__9758 (
            .O(N__39343),
            .I(N__38969));
    ClkMux I__9757 (
            .O(N__39342),
            .I(N__38969));
    ClkMux I__9756 (
            .O(N__39341),
            .I(N__38969));
    ClkMux I__9755 (
            .O(N__39340),
            .I(N__38969));
    ClkMux I__9754 (
            .O(N__39339),
            .I(N__38969));
    ClkMux I__9753 (
            .O(N__39338),
            .I(N__38969));
    ClkMux I__9752 (
            .O(N__39337),
            .I(N__38969));
    ClkMux I__9751 (
            .O(N__39336),
            .I(N__38969));
    ClkMux I__9750 (
            .O(N__39335),
            .I(N__38969));
    ClkMux I__9749 (
            .O(N__39334),
            .I(N__38969));
    ClkMux I__9748 (
            .O(N__39333),
            .I(N__38969));
    ClkMux I__9747 (
            .O(N__39332),
            .I(N__38969));
    ClkMux I__9746 (
            .O(N__39331),
            .I(N__38969));
    ClkMux I__9745 (
            .O(N__39330),
            .I(N__38969));
    ClkMux I__9744 (
            .O(N__39329),
            .I(N__38969));
    ClkMux I__9743 (
            .O(N__39328),
            .I(N__38969));
    ClkMux I__9742 (
            .O(N__39327),
            .I(N__38969));
    ClkMux I__9741 (
            .O(N__39326),
            .I(N__38969));
    ClkMux I__9740 (
            .O(N__39325),
            .I(N__38969));
    ClkMux I__9739 (
            .O(N__39324),
            .I(N__38969));
    ClkMux I__9738 (
            .O(N__39323),
            .I(N__38969));
    ClkMux I__9737 (
            .O(N__39322),
            .I(N__38969));
    ClkMux I__9736 (
            .O(N__39321),
            .I(N__38969));
    ClkMux I__9735 (
            .O(N__39320),
            .I(N__38969));
    ClkMux I__9734 (
            .O(N__39319),
            .I(N__38969));
    ClkMux I__9733 (
            .O(N__39318),
            .I(N__38969));
    ClkMux I__9732 (
            .O(N__39317),
            .I(N__38969));
    ClkMux I__9731 (
            .O(N__39316),
            .I(N__38969));
    ClkMux I__9730 (
            .O(N__39315),
            .I(N__38969));
    ClkMux I__9729 (
            .O(N__39314),
            .I(N__38969));
    ClkMux I__9728 (
            .O(N__39313),
            .I(N__38969));
    ClkMux I__9727 (
            .O(N__39312),
            .I(N__38969));
    ClkMux I__9726 (
            .O(N__39311),
            .I(N__38969));
    ClkMux I__9725 (
            .O(N__39310),
            .I(N__38969));
    ClkMux I__9724 (
            .O(N__39309),
            .I(N__38969));
    ClkMux I__9723 (
            .O(N__39308),
            .I(N__38969));
    ClkMux I__9722 (
            .O(N__39307),
            .I(N__38969));
    ClkMux I__9721 (
            .O(N__39306),
            .I(N__38969));
    ClkMux I__9720 (
            .O(N__39305),
            .I(N__38969));
    ClkMux I__9719 (
            .O(N__39304),
            .I(N__38969));
    ClkMux I__9718 (
            .O(N__39303),
            .I(N__38969));
    ClkMux I__9717 (
            .O(N__39302),
            .I(N__38969));
    ClkMux I__9716 (
            .O(N__39301),
            .I(N__38969));
    ClkMux I__9715 (
            .O(N__39300),
            .I(N__38969));
    ClkMux I__9714 (
            .O(N__39299),
            .I(N__38969));
    ClkMux I__9713 (
            .O(N__39298),
            .I(N__38969));
    ClkMux I__9712 (
            .O(N__39297),
            .I(N__38969));
    ClkMux I__9711 (
            .O(N__39296),
            .I(N__38969));
    ClkMux I__9710 (
            .O(N__39295),
            .I(N__38969));
    ClkMux I__9709 (
            .O(N__39294),
            .I(N__38969));
    ClkMux I__9708 (
            .O(N__39293),
            .I(N__38969));
    ClkMux I__9707 (
            .O(N__39292),
            .I(N__38969));
    ClkMux I__9706 (
            .O(N__39291),
            .I(N__38969));
    ClkMux I__9705 (
            .O(N__39290),
            .I(N__38969));
    ClkMux I__9704 (
            .O(N__39289),
            .I(N__38969));
    ClkMux I__9703 (
            .O(N__39288),
            .I(N__38969));
    ClkMux I__9702 (
            .O(N__39287),
            .I(N__38969));
    ClkMux I__9701 (
            .O(N__39286),
            .I(N__38969));
    ClkMux I__9700 (
            .O(N__39285),
            .I(N__38969));
    ClkMux I__9699 (
            .O(N__39284),
            .I(N__38969));
    ClkMux I__9698 (
            .O(N__39283),
            .I(N__38969));
    ClkMux I__9697 (
            .O(N__39282),
            .I(N__38969));
    ClkMux I__9696 (
            .O(N__39281),
            .I(N__38969));
    ClkMux I__9695 (
            .O(N__39280),
            .I(N__38969));
    GlobalMux I__9694 (
            .O(N__38969),
            .I(N__38966));
    gio2CtrlBuf I__9693 (
            .O(N__38966),
            .I(clk_0_c_g));
    SRMux I__9692 (
            .O(N__38963),
            .I(N__38924));
    SRMux I__9691 (
            .O(N__38962),
            .I(N__38924));
    SRMux I__9690 (
            .O(N__38961),
            .I(N__38924));
    SRMux I__9689 (
            .O(N__38960),
            .I(N__38924));
    SRMux I__9688 (
            .O(N__38959),
            .I(N__38924));
    SRMux I__9687 (
            .O(N__38958),
            .I(N__38924));
    SRMux I__9686 (
            .O(N__38957),
            .I(N__38924));
    SRMux I__9685 (
            .O(N__38956),
            .I(N__38924));
    SRMux I__9684 (
            .O(N__38955),
            .I(N__38924));
    SRMux I__9683 (
            .O(N__38954),
            .I(N__38924));
    SRMux I__9682 (
            .O(N__38953),
            .I(N__38924));
    SRMux I__9681 (
            .O(N__38952),
            .I(N__38924));
    SRMux I__9680 (
            .O(N__38951),
            .I(N__38924));
    GlobalMux I__9679 (
            .O(N__38924),
            .I(N__38921));
    gio2CtrlBuf I__9678 (
            .O(N__38921),
            .I(N_527_g));
    InMux I__9677 (
            .O(N__38918),
            .I(N__38914));
    InMux I__9676 (
            .O(N__38917),
            .I(N__38911));
    LocalMux I__9675 (
            .O(N__38914),
            .I(N__38904));
    LocalMux I__9674 (
            .O(N__38911),
            .I(N__38904));
    InMux I__9673 (
            .O(N__38910),
            .I(N__38900));
    CascadeMux I__9672 (
            .O(N__38909),
            .I(N__38897));
    Span4Mux_v I__9671 (
            .O(N__38904),
            .I(N__38891));
    InMux I__9670 (
            .O(N__38903),
            .I(N__38887));
    LocalMux I__9669 (
            .O(N__38900),
            .I(N__38883));
    InMux I__9668 (
            .O(N__38897),
            .I(N__38880));
    CascadeMux I__9667 (
            .O(N__38896),
            .I(N__38877));
    InMux I__9666 (
            .O(N__38895),
            .I(N__38874));
    InMux I__9665 (
            .O(N__38894),
            .I(N__38871));
    Span4Mux_h I__9664 (
            .O(N__38891),
            .I(N__38868));
    InMux I__9663 (
            .O(N__38890),
            .I(N__38865));
    LocalMux I__9662 (
            .O(N__38887),
            .I(N__38862));
    InMux I__9661 (
            .O(N__38886),
            .I(N__38859));
    Span4Mux_v I__9660 (
            .O(N__38883),
            .I(N__38856));
    LocalMux I__9659 (
            .O(N__38880),
            .I(N__38853));
    InMux I__9658 (
            .O(N__38877),
            .I(N__38850));
    LocalMux I__9657 (
            .O(N__38874),
            .I(N__38845));
    LocalMux I__9656 (
            .O(N__38871),
            .I(N__38845));
    Span4Mux_v I__9655 (
            .O(N__38868),
            .I(N__38842));
    LocalMux I__9654 (
            .O(N__38865),
            .I(N__38839));
    Span4Mux_v I__9653 (
            .O(N__38862),
            .I(N__38836));
    LocalMux I__9652 (
            .O(N__38859),
            .I(N__38833));
    Span4Mux_h I__9651 (
            .O(N__38856),
            .I(N__38828));
    Span4Mux_v I__9650 (
            .O(N__38853),
            .I(N__38828));
    LocalMux I__9649 (
            .O(N__38850),
            .I(N__38825));
    Span12Mux_h I__9648 (
            .O(N__38845),
            .I(N__38822));
    Span4Mux_v I__9647 (
            .O(N__38842),
            .I(N__38817));
    Span4Mux_v I__9646 (
            .O(N__38839),
            .I(N__38817));
    Span4Mux_h I__9645 (
            .O(N__38836),
            .I(N__38812));
    Span4Mux_v I__9644 (
            .O(N__38833),
            .I(N__38812));
    Span4Mux_h I__9643 (
            .O(N__38828),
            .I(N__38807));
    Span4Mux_v I__9642 (
            .O(N__38825),
            .I(N__38807));
    Span12Mux_h I__9641 (
            .O(N__38822),
            .I(N__38804));
    Sp12to4 I__9640 (
            .O(N__38817),
            .I(N__38801));
    Span4Mux_v I__9639 (
            .O(N__38812),
            .I(N__38796));
    Span4Mux_h I__9638 (
            .O(N__38807),
            .I(N__38796));
    Span12Mux_v I__9637 (
            .O(N__38804),
            .I(N__38793));
    Span12Mux_h I__9636 (
            .O(N__38801),
            .I(N__38790));
    Span4Mux_h I__9635 (
            .O(N__38796),
            .I(N__38787));
    Odrv12 I__9634 (
            .O(N__38793),
            .I(port_data_c_5));
    Odrv12 I__9633 (
            .O(N__38790),
            .I(port_data_c_5));
    Odrv4 I__9632 (
            .O(N__38787),
            .I(port_data_c_5));
    InMux I__9631 (
            .O(N__38780),
            .I(N__38777));
    LocalMux I__9630 (
            .O(N__38777),
            .I(M_this_map_ram_write_data_5));
    InMux I__9629 (
            .O(N__38774),
            .I(N__38770));
    CascadeMux I__9628 (
            .O(N__38773),
            .I(N__38765));
    LocalMux I__9627 (
            .O(N__38770),
            .I(N__38762));
    InMux I__9626 (
            .O(N__38769),
            .I(N__38756));
    InMux I__9625 (
            .O(N__38768),
            .I(N__38753));
    InMux I__9624 (
            .O(N__38765),
            .I(N__38750));
    Span4Mux_v I__9623 (
            .O(N__38762),
            .I(N__38747));
    InMux I__9622 (
            .O(N__38761),
            .I(N__38744));
    InMux I__9621 (
            .O(N__38760),
            .I(N__38741));
    InMux I__9620 (
            .O(N__38759),
            .I(N__38738));
    LocalMux I__9619 (
            .O(N__38756),
            .I(N__38734));
    LocalMux I__9618 (
            .O(N__38753),
            .I(N__38731));
    LocalMux I__9617 (
            .O(N__38750),
            .I(N__38726));
    Span4Mux_v I__9616 (
            .O(N__38747),
            .I(N__38723));
    LocalMux I__9615 (
            .O(N__38744),
            .I(N__38720));
    LocalMux I__9614 (
            .O(N__38741),
            .I(N__38715));
    LocalMux I__9613 (
            .O(N__38738),
            .I(N__38715));
    CascadeMux I__9612 (
            .O(N__38737),
            .I(N__38712));
    Span4Mux_h I__9611 (
            .O(N__38734),
            .I(N__38709));
    Span4Mux_h I__9610 (
            .O(N__38731),
            .I(N__38706));
    InMux I__9609 (
            .O(N__38730),
            .I(N__38703));
    InMux I__9608 (
            .O(N__38729),
            .I(N__38700));
    Span4Mux_v I__9607 (
            .O(N__38726),
            .I(N__38697));
    Span4Mux_v I__9606 (
            .O(N__38723),
            .I(N__38694));
    Span4Mux_v I__9605 (
            .O(N__38720),
            .I(N__38689));
    Span4Mux_h I__9604 (
            .O(N__38715),
            .I(N__38689));
    InMux I__9603 (
            .O(N__38712),
            .I(N__38686));
    Sp12to4 I__9602 (
            .O(N__38709),
            .I(N__38681));
    Sp12to4 I__9601 (
            .O(N__38706),
            .I(N__38681));
    LocalMux I__9600 (
            .O(N__38703),
            .I(N__38676));
    LocalMux I__9599 (
            .O(N__38700),
            .I(N__38676));
    Span4Mux_v I__9598 (
            .O(N__38697),
            .I(N__38667));
    Span4Mux_h I__9597 (
            .O(N__38694),
            .I(N__38667));
    Span4Mux_h I__9596 (
            .O(N__38689),
            .I(N__38667));
    LocalMux I__9595 (
            .O(N__38686),
            .I(N__38667));
    Span12Mux_s10_v I__9594 (
            .O(N__38681),
            .I(N__38664));
    Span12Mux_s10_v I__9593 (
            .O(N__38676),
            .I(N__38661));
    Span4Mux_v I__9592 (
            .O(N__38667),
            .I(N__38658));
    Span12Mux_v I__9591 (
            .O(N__38664),
            .I(N__38655));
    Span12Mux_v I__9590 (
            .O(N__38661),
            .I(N__38652));
    Span4Mux_v I__9589 (
            .O(N__38658),
            .I(N__38649));
    Span12Mux_h I__9588 (
            .O(N__38655),
            .I(N__38646));
    Span12Mux_h I__9587 (
            .O(N__38652),
            .I(N__38641));
    Sp12to4 I__9586 (
            .O(N__38649),
            .I(N__38641));
    Odrv12 I__9585 (
            .O(N__38646),
            .I(port_data_c_7));
    Odrv12 I__9584 (
            .O(N__38641),
            .I(port_data_c_7));
    InMux I__9583 (
            .O(N__38636),
            .I(N__38633));
    LocalMux I__9582 (
            .O(N__38633),
            .I(M_this_map_ram_write_data_7));
    CEMux I__9581 (
            .O(N__38630),
            .I(N__38621));
    InMux I__9580 (
            .O(N__38629),
            .I(N__38609));
    InMux I__9579 (
            .O(N__38628),
            .I(N__38609));
    InMux I__9578 (
            .O(N__38627),
            .I(N__38609));
    InMux I__9577 (
            .O(N__38626),
            .I(N__38609));
    CEMux I__9576 (
            .O(N__38625),
            .I(N__38606));
    InMux I__9575 (
            .O(N__38624),
            .I(N__38603));
    LocalMux I__9574 (
            .O(N__38621),
            .I(N__38599));
    InMux I__9573 (
            .O(N__38620),
            .I(N__38596));
    InMux I__9572 (
            .O(N__38619),
            .I(N__38591));
    InMux I__9571 (
            .O(N__38618),
            .I(N__38591));
    LocalMux I__9570 (
            .O(N__38609),
            .I(N__38588));
    LocalMux I__9569 (
            .O(N__38606),
            .I(N__38584));
    LocalMux I__9568 (
            .O(N__38603),
            .I(N__38581));
    CascadeMux I__9567 (
            .O(N__38602),
            .I(N__38578));
    Span4Mux_h I__9566 (
            .O(N__38599),
            .I(N__38573));
    LocalMux I__9565 (
            .O(N__38596),
            .I(N__38573));
    LocalMux I__9564 (
            .O(N__38591),
            .I(N__38570));
    Span4Mux_h I__9563 (
            .O(N__38588),
            .I(N__38567));
    InMux I__9562 (
            .O(N__38587),
            .I(N__38564));
    Span4Mux_v I__9561 (
            .O(N__38584),
            .I(N__38559));
    Span4Mux_h I__9560 (
            .O(N__38581),
            .I(N__38559));
    InMux I__9559 (
            .O(N__38578),
            .I(N__38556));
    Span4Mux_v I__9558 (
            .O(N__38573),
            .I(N__38553));
    Span4Mux_v I__9557 (
            .O(N__38570),
            .I(N__38550));
    Span4Mux_v I__9556 (
            .O(N__38567),
            .I(N__38547));
    LocalMux I__9555 (
            .O(N__38564),
            .I(N__38540));
    Sp12to4 I__9554 (
            .O(N__38559),
            .I(N__38540));
    LocalMux I__9553 (
            .O(N__38556),
            .I(N__38540));
    Span4Mux_h I__9552 (
            .O(N__38553),
            .I(N__38537));
    Sp12to4 I__9551 (
            .O(N__38550),
            .I(N__38530));
    Sp12to4 I__9550 (
            .O(N__38547),
            .I(N__38530));
    Span12Mux_v I__9549 (
            .O(N__38540),
            .I(N__38530));
    Span4Mux_h I__9548 (
            .O(N__38537),
            .I(N__38527));
    Span12Mux_h I__9547 (
            .O(N__38530),
            .I(N__38524));
    Odrv4 I__9546 (
            .O(N__38527),
            .I(M_this_state_d_0_sqmuxa));
    Odrv12 I__9545 (
            .O(N__38524),
            .I(M_this_state_d_0_sqmuxa));
    CascadeMux I__9544 (
            .O(N__38519),
            .I(N__38516));
    CascadeBuf I__9543 (
            .O(N__38516),
            .I(N__38513));
    CascadeMux I__9542 (
            .O(N__38513),
            .I(N__38510));
    InMux I__9541 (
            .O(N__38510),
            .I(N__38506));
    InMux I__9540 (
            .O(N__38509),
            .I(N__38503));
    LocalMux I__9539 (
            .O(N__38506),
            .I(N__38500));
    LocalMux I__9538 (
            .O(N__38503),
            .I(N__38495));
    Span4Mux_v I__9537 (
            .O(N__38500),
            .I(N__38495));
    Odrv4 I__9536 (
            .O(N__38495),
            .I(M_this_map_address_qZ0Z_0));
    CascadeMux I__9535 (
            .O(N__38492),
            .I(N__38489));
    CascadeBuf I__9534 (
            .O(N__38489),
            .I(N__38486));
    CascadeMux I__9533 (
            .O(N__38486),
            .I(N__38483));
    InMux I__9532 (
            .O(N__38483),
            .I(N__38480));
    LocalMux I__9531 (
            .O(N__38480),
            .I(N__38476));
    InMux I__9530 (
            .O(N__38479),
            .I(N__38473));
    Span4Mux_v I__9529 (
            .O(N__38476),
            .I(N__38470));
    LocalMux I__9528 (
            .O(N__38473),
            .I(M_this_map_address_qZ0Z_1));
    Odrv4 I__9527 (
            .O(N__38470),
            .I(M_this_map_address_qZ0Z_1));
    InMux I__9526 (
            .O(N__38465),
            .I(un1_M_this_map_address_q_cry_0));
    CascadeMux I__9525 (
            .O(N__38462),
            .I(N__38459));
    CascadeBuf I__9524 (
            .O(N__38459),
            .I(N__38456));
    CascadeMux I__9523 (
            .O(N__38456),
            .I(N__38453));
    InMux I__9522 (
            .O(N__38453),
            .I(N__38450));
    LocalMux I__9521 (
            .O(N__38450),
            .I(N__38446));
    InMux I__9520 (
            .O(N__38449),
            .I(N__38443));
    Span4Mux_h I__9519 (
            .O(N__38446),
            .I(N__38440));
    LocalMux I__9518 (
            .O(N__38443),
            .I(M_this_map_address_qZ0Z_2));
    Odrv4 I__9517 (
            .O(N__38440),
            .I(M_this_map_address_qZ0Z_2));
    InMux I__9516 (
            .O(N__38435),
            .I(un1_M_this_map_address_q_cry_1));
    CascadeMux I__9515 (
            .O(N__38432),
            .I(N__38429));
    CascadeBuf I__9514 (
            .O(N__38429),
            .I(N__38426));
    CascadeMux I__9513 (
            .O(N__38426),
            .I(N__38423));
    InMux I__9512 (
            .O(N__38423),
            .I(N__38419));
    InMux I__9511 (
            .O(N__38422),
            .I(N__38416));
    LocalMux I__9510 (
            .O(N__38419),
            .I(N__38413));
    LocalMux I__9509 (
            .O(N__38416),
            .I(M_this_map_address_qZ0Z_3));
    Odrv4 I__9508 (
            .O(N__38413),
            .I(M_this_map_address_qZ0Z_3));
    InMux I__9507 (
            .O(N__38408),
            .I(un1_M_this_map_address_q_cry_2));
    CascadeMux I__9506 (
            .O(N__38405),
            .I(N__38402));
    CascadeBuf I__9505 (
            .O(N__38402),
            .I(N__38399));
    CascadeMux I__9504 (
            .O(N__38399),
            .I(N__38396));
    InMux I__9503 (
            .O(N__38396),
            .I(N__38393));
    LocalMux I__9502 (
            .O(N__38393),
            .I(N__38389));
    InMux I__9501 (
            .O(N__38392),
            .I(N__38386));
    Span4Mux_h I__9500 (
            .O(N__38389),
            .I(N__38383));
    LocalMux I__9499 (
            .O(N__38386),
            .I(M_this_map_address_qZ0Z_4));
    Odrv4 I__9498 (
            .O(N__38383),
            .I(M_this_map_address_qZ0Z_4));
    InMux I__9497 (
            .O(N__38378),
            .I(un1_M_this_map_address_q_cry_3));
    CascadeMux I__9496 (
            .O(N__38375),
            .I(N__38372));
    CascadeBuf I__9495 (
            .O(N__38372),
            .I(N__38369));
    CascadeMux I__9494 (
            .O(N__38369),
            .I(N__38366));
    InMux I__9493 (
            .O(N__38366),
            .I(N__38362));
    InMux I__9492 (
            .O(N__38365),
            .I(N__38359));
    LocalMux I__9491 (
            .O(N__38362),
            .I(N__38356));
    LocalMux I__9490 (
            .O(N__38359),
            .I(M_this_map_address_qZ0Z_5));
    Odrv4 I__9489 (
            .O(N__38356),
            .I(M_this_map_address_qZ0Z_5));
    InMux I__9488 (
            .O(N__38351),
            .I(un1_M_this_map_address_q_cry_4));
    InMux I__9487 (
            .O(N__38348),
            .I(N__38340));
    InMux I__9486 (
            .O(N__38347),
            .I(N__38335));
    InMux I__9485 (
            .O(N__38346),
            .I(N__38335));
    InMux I__9484 (
            .O(N__38345),
            .I(N__38329));
    InMux I__9483 (
            .O(N__38344),
            .I(N__38329));
    InMux I__9482 (
            .O(N__38343),
            .I(N__38326));
    LocalMux I__9481 (
            .O(N__38340),
            .I(N__38323));
    LocalMux I__9480 (
            .O(N__38335),
            .I(N__38320));
    InMux I__9479 (
            .O(N__38334),
            .I(N__38317));
    LocalMux I__9478 (
            .O(N__38329),
            .I(N__38312));
    LocalMux I__9477 (
            .O(N__38326),
            .I(N__38312));
    Span4Mux_h I__9476 (
            .O(N__38323),
            .I(N__38309));
    Span4Mux_v I__9475 (
            .O(N__38320),
            .I(N__38301));
    LocalMux I__9474 (
            .O(N__38317),
            .I(N__38301));
    Span4Mux_v I__9473 (
            .O(N__38312),
            .I(N__38301));
    Span4Mux_v I__9472 (
            .O(N__38309),
            .I(N__38298));
    InMux I__9471 (
            .O(N__38308),
            .I(N__38295));
    Span4Mux_h I__9470 (
            .O(N__38301),
            .I(N__38292));
    Odrv4 I__9469 (
            .O(N__38298),
            .I(N_930));
    LocalMux I__9468 (
            .O(N__38295),
            .I(N_930));
    Odrv4 I__9467 (
            .O(N__38292),
            .I(N_930));
    InMux I__9466 (
            .O(N__38285),
            .I(N__38274));
    InMux I__9465 (
            .O(N__38284),
            .I(N__38271));
    InMux I__9464 (
            .O(N__38283),
            .I(N__38268));
    InMux I__9463 (
            .O(N__38282),
            .I(N__38264));
    InMux I__9462 (
            .O(N__38281),
            .I(N__38261));
    InMux I__9461 (
            .O(N__38280),
            .I(N__38258));
    InMux I__9460 (
            .O(N__38279),
            .I(N__38255));
    InMux I__9459 (
            .O(N__38278),
            .I(N__38252));
    InMux I__9458 (
            .O(N__38277),
            .I(N__38249));
    LocalMux I__9457 (
            .O(N__38274),
            .I(N__38244));
    LocalMux I__9456 (
            .O(N__38271),
            .I(N__38244));
    LocalMux I__9455 (
            .O(N__38268),
            .I(N__38241));
    InMux I__9454 (
            .O(N__38267),
            .I(N__38238));
    LocalMux I__9453 (
            .O(N__38264),
            .I(N__38235));
    LocalMux I__9452 (
            .O(N__38261),
            .I(N__38230));
    LocalMux I__9451 (
            .O(N__38258),
            .I(N__38230));
    LocalMux I__9450 (
            .O(N__38255),
            .I(N__38222));
    LocalMux I__9449 (
            .O(N__38252),
            .I(N__38222));
    LocalMux I__9448 (
            .O(N__38249),
            .I(N__38219));
    Span4Mux_v I__9447 (
            .O(N__38244),
            .I(N__38214));
    Span4Mux_v I__9446 (
            .O(N__38241),
            .I(N__38214));
    LocalMux I__9445 (
            .O(N__38238),
            .I(N__38211));
    Span4Mux_v I__9444 (
            .O(N__38235),
            .I(N__38206));
    Span4Mux_h I__9443 (
            .O(N__38230),
            .I(N__38206));
    InMux I__9442 (
            .O(N__38229),
            .I(N__38203));
    InMux I__9441 (
            .O(N__38228),
            .I(N__38198));
    InMux I__9440 (
            .O(N__38227),
            .I(N__38198));
    Span12Mux_h I__9439 (
            .O(N__38222),
            .I(N__38195));
    Span4Mux_v I__9438 (
            .O(N__38219),
            .I(N__38192));
    Span4Mux_h I__9437 (
            .O(N__38214),
            .I(N__38185));
    Span4Mux_v I__9436 (
            .O(N__38211),
            .I(N__38185));
    Span4Mux_v I__9435 (
            .O(N__38206),
            .I(N__38185));
    LocalMux I__9434 (
            .O(N__38203),
            .I(N__38180));
    LocalMux I__9433 (
            .O(N__38198),
            .I(N__38180));
    Odrv12 I__9432 (
            .O(N__38195),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__9431 (
            .O(N__38192),
            .I(M_this_state_qZ0Z_9));
    Odrv4 I__9430 (
            .O(N__38185),
            .I(M_this_state_qZ0Z_9));
    Odrv12 I__9429 (
            .O(N__38180),
            .I(M_this_state_qZ0Z_9));
    InMux I__9428 (
            .O(N__38171),
            .I(N__38168));
    LocalMux I__9427 (
            .O(N__38168),
            .I(N__38165));
    Span4Mux_h I__9426 (
            .O(N__38165),
            .I(N__38161));
    InMux I__9425 (
            .O(N__38164),
            .I(N__38156));
    Span4Mux_h I__9424 (
            .O(N__38161),
            .I(N__38153));
    InMux I__9423 (
            .O(N__38160),
            .I(N__38148));
    InMux I__9422 (
            .O(N__38159),
            .I(N__38148));
    LocalMux I__9421 (
            .O(N__38156),
            .I(M_this_state_qZ0Z_4));
    Odrv4 I__9420 (
            .O(N__38153),
            .I(M_this_state_qZ0Z_4));
    LocalMux I__9419 (
            .O(N__38148),
            .I(M_this_state_qZ0Z_4));
    CascadeMux I__9418 (
            .O(N__38141),
            .I(N__38138));
    InMux I__9417 (
            .O(N__38138),
            .I(N__38135));
    LocalMux I__9416 (
            .O(N__38135),
            .I(N__38132));
    Odrv4 I__9415 (
            .O(N__38132),
            .I(\this_start_data_delay.N_332 ));
    InMux I__9414 (
            .O(N__38129),
            .I(N__38124));
    InMux I__9413 (
            .O(N__38128),
            .I(N__38121));
    InMux I__9412 (
            .O(N__38127),
            .I(N__38118));
    LocalMux I__9411 (
            .O(N__38124),
            .I(N__38113));
    LocalMux I__9410 (
            .O(N__38121),
            .I(N__38110));
    LocalMux I__9409 (
            .O(N__38118),
            .I(N__38107));
    InMux I__9408 (
            .O(N__38117),
            .I(N__38104));
    InMux I__9407 (
            .O(N__38116),
            .I(N__38098));
    Span4Mux_h I__9406 (
            .O(N__38113),
            .I(N__38093));
    Span4Mux_h I__9405 (
            .O(N__38110),
            .I(N__38093));
    Span4Mux_h I__9404 (
            .O(N__38107),
            .I(N__38088));
    LocalMux I__9403 (
            .O(N__38104),
            .I(N__38088));
    InMux I__9402 (
            .O(N__38103),
            .I(N__38085));
    InMux I__9401 (
            .O(N__38102),
            .I(N__38082));
    InMux I__9400 (
            .O(N__38101),
            .I(N__38079));
    LocalMux I__9399 (
            .O(N__38098),
            .I(N__38075));
    Span4Mux_v I__9398 (
            .O(N__38093),
            .I(N__38072));
    Span4Mux_h I__9397 (
            .O(N__38088),
            .I(N__38069));
    LocalMux I__9396 (
            .O(N__38085),
            .I(N__38066));
    LocalMux I__9395 (
            .O(N__38082),
            .I(N__38061));
    LocalMux I__9394 (
            .O(N__38079),
            .I(N__38061));
    InMux I__9393 (
            .O(N__38078),
            .I(N__38058));
    Span12Mux_h I__9392 (
            .O(N__38075),
            .I(N__38055));
    Span4Mux_v I__9391 (
            .O(N__38072),
            .I(N__38052));
    Span4Mux_v I__9390 (
            .O(N__38069),
            .I(N__38049));
    Span4Mux_v I__9389 (
            .O(N__38066),
            .I(N__38042));
    Span4Mux_s3_v I__9388 (
            .O(N__38061),
            .I(N__38042));
    LocalMux I__9387 (
            .O(N__38058),
            .I(N__38042));
    Span12Mux_v I__9386 (
            .O(N__38055),
            .I(N__38039));
    Span4Mux_v I__9385 (
            .O(N__38052),
            .I(N__38036));
    Span4Mux_h I__9384 (
            .O(N__38049),
            .I(N__38031));
    Span4Mux_h I__9383 (
            .O(N__38042),
            .I(N__38031));
    Odrv12 I__9382 (
            .O(N__38039),
            .I(port_data_c_0));
    Odrv4 I__9381 (
            .O(N__38036),
            .I(port_data_c_0));
    Odrv4 I__9380 (
            .O(N__38031),
            .I(port_data_c_0));
    InMux I__9379 (
            .O(N__38024),
            .I(N__38021));
    LocalMux I__9378 (
            .O(N__38021),
            .I(N__38018));
    Span4Mux_h I__9377 (
            .O(N__38018),
            .I(N__38015));
    Odrv4 I__9376 (
            .O(N__38015),
            .I(M_this_map_ram_write_data_0));
    IoInMux I__9375 (
            .O(N__38012),
            .I(N__38009));
    LocalMux I__9374 (
            .O(N__38009),
            .I(N__38004));
    InMux I__9373 (
            .O(N__38008),
            .I(N__38001));
    InMux I__9372 (
            .O(N__38007),
            .I(N__37998));
    Span12Mux_s11_h I__9371 (
            .O(N__38004),
            .I(N__37993));
    LocalMux I__9370 (
            .O(N__38001),
            .I(N__37990));
    LocalMux I__9369 (
            .O(N__37998),
            .I(N__37987));
    InMux I__9368 (
            .O(N__37997),
            .I(N__37984));
    CascadeMux I__9367 (
            .O(N__37996),
            .I(N__37980));
    Span12Mux_v I__9366 (
            .O(N__37993),
            .I(N__37975));
    Span12Mux_v I__9365 (
            .O(N__37990),
            .I(N__37972));
    Span4Mux_h I__9364 (
            .O(N__37987),
            .I(N__37969));
    LocalMux I__9363 (
            .O(N__37984),
            .I(N__37966));
    InMux I__9362 (
            .O(N__37983),
            .I(N__37961));
    InMux I__9361 (
            .O(N__37980),
            .I(N__37961));
    InMux I__9360 (
            .O(N__37979),
            .I(N__37956));
    InMux I__9359 (
            .O(N__37978),
            .I(N__37956));
    Odrv12 I__9358 (
            .O(N__37975),
            .I(led_c_1));
    Odrv12 I__9357 (
            .O(N__37972),
            .I(led_c_1));
    Odrv4 I__9356 (
            .O(N__37969),
            .I(led_c_1));
    Odrv4 I__9355 (
            .O(N__37966),
            .I(led_c_1));
    LocalMux I__9354 (
            .O(N__37961),
            .I(led_c_1));
    LocalMux I__9353 (
            .O(N__37956),
            .I(led_c_1));
    InMux I__9352 (
            .O(N__37943),
            .I(N__37940));
    LocalMux I__9351 (
            .O(N__37940),
            .I(N__37935));
    InMux I__9350 (
            .O(N__37939),
            .I(N__37932));
    CascadeMux I__9349 (
            .O(N__37938),
            .I(N__37929));
    Span4Mux_h I__9348 (
            .O(N__37935),
            .I(N__37926));
    LocalMux I__9347 (
            .O(N__37932),
            .I(N__37923));
    InMux I__9346 (
            .O(N__37929),
            .I(N__37920));
    Odrv4 I__9345 (
            .O(N__37926),
            .I(N_466));
    Odrv12 I__9344 (
            .O(N__37923),
            .I(N_466));
    LocalMux I__9343 (
            .O(N__37920),
            .I(N_466));
    IoInMux I__9342 (
            .O(N__37913),
            .I(N__37910));
    LocalMux I__9341 (
            .O(N__37910),
            .I(N__37907));
    Span12Mux_s9_h I__9340 (
            .O(N__37907),
            .I(N__37904));
    Span12Mux_v I__9339 (
            .O(N__37904),
            .I(N__37901));
    Odrv12 I__9338 (
            .O(N__37901),
            .I(led_c_7));
    InMux I__9337 (
            .O(N__37898),
            .I(N__37895));
    LocalMux I__9336 (
            .O(N__37895),
            .I(N__37892));
    Span4Mux_v I__9335 (
            .O(N__37892),
            .I(N__37888));
    InMux I__9334 (
            .O(N__37891),
            .I(N__37885));
    Span4Mux_h I__9333 (
            .O(N__37888),
            .I(N__37880));
    LocalMux I__9332 (
            .O(N__37885),
            .I(N__37880));
    Span4Mux_h I__9331 (
            .O(N__37880),
            .I(N__37875));
    InMux I__9330 (
            .O(N__37879),
            .I(N__37871));
    InMux I__9329 (
            .O(N__37878),
            .I(N__37868));
    Span4Mux_v I__9328 (
            .O(N__37875),
            .I(N__37865));
    InMux I__9327 (
            .O(N__37874),
            .I(N__37862));
    LocalMux I__9326 (
            .O(N__37871),
            .I(N__37857));
    LocalMux I__9325 (
            .O(N__37868),
            .I(N__37854));
    Span4Mux_v I__9324 (
            .O(N__37865),
            .I(N__37847));
    LocalMux I__9323 (
            .O(N__37862),
            .I(N__37847));
    InMux I__9322 (
            .O(N__37861),
            .I(N__37844));
    InMux I__9321 (
            .O(N__37860),
            .I(N__37841));
    Span4Mux_v I__9320 (
            .O(N__37857),
            .I(N__37838));
    Span4Mux_v I__9319 (
            .O(N__37854),
            .I(N__37835));
    InMux I__9318 (
            .O(N__37853),
            .I(N__37832));
    InMux I__9317 (
            .O(N__37852),
            .I(N__37829));
    Span4Mux_v I__9316 (
            .O(N__37847),
            .I(N__37826));
    LocalMux I__9315 (
            .O(N__37844),
            .I(N__37823));
    LocalMux I__9314 (
            .O(N__37841),
            .I(N__37820));
    Sp12to4 I__9313 (
            .O(N__37838),
            .I(N__37817));
    Span4Mux_h I__9312 (
            .O(N__37835),
            .I(N__37814));
    LocalMux I__9311 (
            .O(N__37832),
            .I(N__37809));
    LocalMux I__9310 (
            .O(N__37829),
            .I(N__37809));
    Span4Mux_h I__9309 (
            .O(N__37826),
            .I(N__37804));
    Span4Mux_v I__9308 (
            .O(N__37823),
            .I(N__37804));
    Span12Mux_h I__9307 (
            .O(N__37820),
            .I(N__37801));
    Span12Mux_h I__9306 (
            .O(N__37817),
            .I(N__37798));
    Sp12to4 I__9305 (
            .O(N__37814),
            .I(N__37793));
    Span12Mux_h I__9304 (
            .O(N__37809),
            .I(N__37793));
    Span4Mux_v I__9303 (
            .O(N__37804),
            .I(N__37790));
    Span12Mux_h I__9302 (
            .O(N__37801),
            .I(N__37787));
    Span12Mux_v I__9301 (
            .O(N__37798),
            .I(N__37782));
    Span12Mux_h I__9300 (
            .O(N__37793),
            .I(N__37782));
    Span4Mux_h I__9299 (
            .O(N__37790),
            .I(N__37779));
    Odrv12 I__9298 (
            .O(N__37787),
            .I(port_data_c_3));
    Odrv12 I__9297 (
            .O(N__37782),
            .I(port_data_c_3));
    Odrv4 I__9296 (
            .O(N__37779),
            .I(port_data_c_3));
    InMux I__9295 (
            .O(N__37772),
            .I(N__37769));
    LocalMux I__9294 (
            .O(N__37769),
            .I(M_this_map_ram_write_data_3));
    InMux I__9293 (
            .O(N__37766),
            .I(N__37763));
    LocalMux I__9292 (
            .O(N__37763),
            .I(N__37760));
    Span4Mux_v I__9291 (
            .O(N__37760),
            .I(N__37756));
    InMux I__9290 (
            .O(N__37759),
            .I(N__37753));
    Span4Mux_h I__9289 (
            .O(N__37756),
            .I(N__37746));
    LocalMux I__9288 (
            .O(N__37753),
            .I(N__37746));
    InMux I__9287 (
            .O(N__37752),
            .I(N__37743));
    InMux I__9286 (
            .O(N__37751),
            .I(N__37740));
    Span4Mux_h I__9285 (
            .O(N__37746),
            .I(N__37736));
    LocalMux I__9284 (
            .O(N__37743),
            .I(N__37731));
    LocalMux I__9283 (
            .O(N__37740),
            .I(N__37728));
    InMux I__9282 (
            .O(N__37739),
            .I(N__37725));
    Span4Mux_v I__9281 (
            .O(N__37736),
            .I(N__37722));
    InMux I__9280 (
            .O(N__37735),
            .I(N__37719));
    InMux I__9279 (
            .O(N__37734),
            .I(N__37716));
    Span4Mux_v I__9278 (
            .O(N__37731),
            .I(N__37712));
    Span4Mux_v I__9277 (
            .O(N__37728),
            .I(N__37709));
    LocalMux I__9276 (
            .O(N__37725),
            .I(N__37706));
    Span4Mux_v I__9275 (
            .O(N__37722),
            .I(N__37701));
    LocalMux I__9274 (
            .O(N__37719),
            .I(N__37701));
    LocalMux I__9273 (
            .O(N__37716),
            .I(N__37698));
    InMux I__9272 (
            .O(N__37715),
            .I(N__37695));
    Sp12to4 I__9271 (
            .O(N__37712),
            .I(N__37689));
    Sp12to4 I__9270 (
            .O(N__37709),
            .I(N__37689));
    Span4Mux_v I__9269 (
            .O(N__37706),
            .I(N__37686));
    Span4Mux_v I__9268 (
            .O(N__37701),
            .I(N__37679));
    Span4Mux_h I__9267 (
            .O(N__37698),
            .I(N__37679));
    LocalMux I__9266 (
            .O(N__37695),
            .I(N__37679));
    InMux I__9265 (
            .O(N__37694),
            .I(N__37676));
    Span12Mux_h I__9264 (
            .O(N__37689),
            .I(N__37671));
    Sp12to4 I__9263 (
            .O(N__37686),
            .I(N__37671));
    IoSpan4Mux I__9262 (
            .O(N__37679),
            .I(N__37668));
    LocalMux I__9261 (
            .O(N__37676),
            .I(N__37665));
    Odrv12 I__9260 (
            .O(N__37671),
            .I(port_data_c_1));
    Odrv4 I__9259 (
            .O(N__37668),
            .I(port_data_c_1));
    Odrv12 I__9258 (
            .O(N__37665),
            .I(port_data_c_1));
    InMux I__9257 (
            .O(N__37658),
            .I(N__37655));
    LocalMux I__9256 (
            .O(N__37655),
            .I(M_this_map_ram_write_data_1));
    InMux I__9255 (
            .O(N__37652),
            .I(N__37646));
    InMux I__9254 (
            .O(N__37651),
            .I(N__37643));
    InMux I__9253 (
            .O(N__37650),
            .I(N__37640));
    InMux I__9252 (
            .O(N__37649),
            .I(N__37637));
    LocalMux I__9251 (
            .O(N__37646),
            .I(N__37634));
    LocalMux I__9250 (
            .O(N__37643),
            .I(N__37629));
    LocalMux I__9249 (
            .O(N__37640),
            .I(N__37625));
    LocalMux I__9248 (
            .O(N__37637),
            .I(N__37622));
    Span4Mux_v I__9247 (
            .O(N__37634),
            .I(N__37619));
    InMux I__9246 (
            .O(N__37633),
            .I(N__37616));
    InMux I__9245 (
            .O(N__37632),
            .I(N__37612));
    Span4Mux_h I__9244 (
            .O(N__37629),
            .I(N__37608));
    InMux I__9243 (
            .O(N__37628),
            .I(N__37605));
    Span4Mux_v I__9242 (
            .O(N__37625),
            .I(N__37602));
    Span4Mux_v I__9241 (
            .O(N__37622),
            .I(N__37599));
    Span4Mux_v I__9240 (
            .O(N__37619),
            .I(N__37594));
    LocalMux I__9239 (
            .O(N__37616),
            .I(N__37594));
    InMux I__9238 (
            .O(N__37615),
            .I(N__37591));
    LocalMux I__9237 (
            .O(N__37612),
            .I(N__37588));
    InMux I__9236 (
            .O(N__37611),
            .I(N__37585));
    Span4Mux_h I__9235 (
            .O(N__37608),
            .I(N__37582));
    LocalMux I__9234 (
            .O(N__37605),
            .I(N__37579));
    Span4Mux_h I__9233 (
            .O(N__37602),
            .I(N__37576));
    Span4Mux_h I__9232 (
            .O(N__37599),
            .I(N__37571));
    Span4Mux_v I__9231 (
            .O(N__37594),
            .I(N__37571));
    LocalMux I__9230 (
            .O(N__37591),
            .I(N__37568));
    Span4Mux_h I__9229 (
            .O(N__37588),
            .I(N__37563));
    LocalMux I__9228 (
            .O(N__37585),
            .I(N__37563));
    Sp12to4 I__9227 (
            .O(N__37582),
            .I(N__37560));
    Span12Mux_v I__9226 (
            .O(N__37579),
            .I(N__37551));
    Sp12to4 I__9225 (
            .O(N__37576),
            .I(N__37551));
    Sp12to4 I__9224 (
            .O(N__37571),
            .I(N__37551));
    Span12Mux_h I__9223 (
            .O(N__37568),
            .I(N__37551));
    Span4Mux_h I__9222 (
            .O(N__37563),
            .I(N__37548));
    Span12Mux_v I__9221 (
            .O(N__37560),
            .I(N__37543));
    Span12Mux_h I__9220 (
            .O(N__37551),
            .I(N__37543));
    Span4Mux_v I__9219 (
            .O(N__37548),
            .I(N__37540));
    Odrv12 I__9218 (
            .O(N__37543),
            .I(port_data_c_2));
    Odrv4 I__9217 (
            .O(N__37540),
            .I(port_data_c_2));
    InMux I__9216 (
            .O(N__37535),
            .I(N__37532));
    LocalMux I__9215 (
            .O(N__37532),
            .I(M_this_map_ram_write_data_2));
    InMux I__9214 (
            .O(N__37529),
            .I(N__37526));
    LocalMux I__9213 (
            .O(N__37526),
            .I(N__37523));
    Span4Mux_v I__9212 (
            .O(N__37523),
            .I(N__37517));
    InMux I__9211 (
            .O(N__37522),
            .I(N__37514));
    CascadeMux I__9210 (
            .O(N__37521),
            .I(N__37511));
    InMux I__9209 (
            .O(N__37520),
            .I(N__37508));
    Span4Mux_v I__9208 (
            .O(N__37517),
            .I(N__37503));
    LocalMux I__9207 (
            .O(N__37514),
            .I(N__37500));
    InMux I__9206 (
            .O(N__37511),
            .I(N__37496));
    LocalMux I__9205 (
            .O(N__37508),
            .I(N__37493));
    InMux I__9204 (
            .O(N__37507),
            .I(N__37490));
    InMux I__9203 (
            .O(N__37506),
            .I(N__37487));
    Span4Mux_v I__9202 (
            .O(N__37503),
            .I(N__37482));
    Span4Mux_v I__9201 (
            .O(N__37500),
            .I(N__37482));
    InMux I__9200 (
            .O(N__37499),
            .I(N__37479));
    LocalMux I__9199 (
            .O(N__37496),
            .I(N__37476));
    Span4Mux_v I__9198 (
            .O(N__37493),
            .I(N__37472));
    LocalMux I__9197 (
            .O(N__37490),
            .I(N__37467));
    LocalMux I__9196 (
            .O(N__37487),
            .I(N__37467));
    Span4Mux_h I__9195 (
            .O(N__37482),
            .I(N__37463));
    LocalMux I__9194 (
            .O(N__37479),
            .I(N__37460));
    Span4Mux_h I__9193 (
            .O(N__37476),
            .I(N__37457));
    InMux I__9192 (
            .O(N__37475),
            .I(N__37454));
    Sp12to4 I__9191 (
            .O(N__37472),
            .I(N__37451));
    Span4Mux_v I__9190 (
            .O(N__37467),
            .I(N__37448));
    InMux I__9189 (
            .O(N__37466),
            .I(N__37445));
    Span4Mux_h I__9188 (
            .O(N__37463),
            .I(N__37440));
    Span4Mux_v I__9187 (
            .O(N__37460),
            .I(N__37440));
    Span4Mux_v I__9186 (
            .O(N__37457),
            .I(N__37435));
    LocalMux I__9185 (
            .O(N__37454),
            .I(N__37435));
    Span12Mux_h I__9184 (
            .O(N__37451),
            .I(N__37432));
    Sp12to4 I__9183 (
            .O(N__37448),
            .I(N__37427));
    LocalMux I__9182 (
            .O(N__37445),
            .I(N__37427));
    Span4Mux_h I__9181 (
            .O(N__37440),
            .I(N__37422));
    Span4Mux_v I__9180 (
            .O(N__37435),
            .I(N__37422));
    Span12Mux_v I__9179 (
            .O(N__37432),
            .I(N__37419));
    Span12Mux_h I__9178 (
            .O(N__37427),
            .I(N__37416));
    Span4Mux_h I__9177 (
            .O(N__37422),
            .I(N__37413));
    Odrv12 I__9176 (
            .O(N__37419),
            .I(port_data_c_4));
    Odrv12 I__9175 (
            .O(N__37416),
            .I(port_data_c_4));
    Odrv4 I__9174 (
            .O(N__37413),
            .I(port_data_c_4));
    InMux I__9173 (
            .O(N__37406),
            .I(N__37403));
    LocalMux I__9172 (
            .O(N__37403),
            .I(N__37400));
    Odrv4 I__9171 (
            .O(N__37400),
            .I(M_this_map_ram_write_data_4));
    InMux I__9170 (
            .O(N__37397),
            .I(N__37393));
    InMux I__9169 (
            .O(N__37396),
            .I(N__37390));
    LocalMux I__9168 (
            .O(N__37393),
            .I(N__37385));
    LocalMux I__9167 (
            .O(N__37390),
            .I(N__37382));
    InMux I__9166 (
            .O(N__37389),
            .I(N__37379));
    InMux I__9165 (
            .O(N__37388),
            .I(N__37376));
    Span4Mux_v I__9164 (
            .O(N__37385),
            .I(N__37368));
    Span4Mux_v I__9163 (
            .O(N__37382),
            .I(N__37368));
    LocalMux I__9162 (
            .O(N__37379),
            .I(N__37368));
    LocalMux I__9161 (
            .O(N__37376),
            .I(N__37365));
    CascadeMux I__9160 (
            .O(N__37375),
            .I(N__37362));
    Span4Mux_v I__9159 (
            .O(N__37368),
            .I(N__37359));
    Span4Mux_h I__9158 (
            .O(N__37365),
            .I(N__37356));
    InMux I__9157 (
            .O(N__37362),
            .I(N__37353));
    Span4Mux_h I__9156 (
            .O(N__37359),
            .I(N__37344));
    Span4Mux_v I__9155 (
            .O(N__37356),
            .I(N__37344));
    LocalMux I__9154 (
            .O(N__37353),
            .I(N__37344));
    InMux I__9153 (
            .O(N__37352),
            .I(N__37341));
    InMux I__9152 (
            .O(N__37351),
            .I(N__37337));
    Span4Mux_v I__9151 (
            .O(N__37344),
            .I(N__37332));
    LocalMux I__9150 (
            .O(N__37341),
            .I(N__37332));
    InMux I__9149 (
            .O(N__37340),
            .I(N__37328));
    LocalMux I__9148 (
            .O(N__37337),
            .I(N__37325));
    Span4Mux_v I__9147 (
            .O(N__37332),
            .I(N__37322));
    CascadeMux I__9146 (
            .O(N__37331),
            .I(N__37319));
    LocalMux I__9145 (
            .O(N__37328),
            .I(N__37316));
    Span4Mux_v I__9144 (
            .O(N__37325),
            .I(N__37313));
    Span4Mux_h I__9143 (
            .O(N__37322),
            .I(N__37309));
    InMux I__9142 (
            .O(N__37319),
            .I(N__37306));
    Span4Mux_h I__9141 (
            .O(N__37316),
            .I(N__37303));
    Span4Mux_h I__9140 (
            .O(N__37313),
            .I(N__37300));
    InMux I__9139 (
            .O(N__37312),
            .I(N__37297));
    Span4Mux_h I__9138 (
            .O(N__37309),
            .I(N__37292));
    LocalMux I__9137 (
            .O(N__37306),
            .I(N__37292));
    Span4Mux_v I__9136 (
            .O(N__37303),
            .I(N__37289));
    Span4Mux_h I__9135 (
            .O(N__37300),
            .I(N__37286));
    LocalMux I__9134 (
            .O(N__37297),
            .I(N__37283));
    Span4Mux_v I__9133 (
            .O(N__37292),
            .I(N__37280));
    Sp12to4 I__9132 (
            .O(N__37289),
            .I(N__37273));
    Sp12to4 I__9131 (
            .O(N__37286),
            .I(N__37273));
    Span12Mux_s9_v I__9130 (
            .O(N__37283),
            .I(N__37273));
    Span4Mux_h I__9129 (
            .O(N__37280),
            .I(N__37270));
    Span12Mux_v I__9128 (
            .O(N__37273),
            .I(N__37267));
    Span4Mux_h I__9127 (
            .O(N__37270),
            .I(N__37264));
    Odrv12 I__9126 (
            .O(N__37267),
            .I(port_data_c_6));
    Odrv4 I__9125 (
            .O(N__37264),
            .I(port_data_c_6));
    InMux I__9124 (
            .O(N__37259),
            .I(N__37256));
    LocalMux I__9123 (
            .O(N__37256),
            .I(N__37253));
    Odrv4 I__9122 (
            .O(N__37253),
            .I(M_this_map_ram_write_data_6));
    IoInMux I__9121 (
            .O(N__37250),
            .I(N__37247));
    LocalMux I__9120 (
            .O(N__37247),
            .I(N__37244));
    Span4Mux_s3_v I__9119 (
            .O(N__37244),
            .I(N__37240));
    CascadeMux I__9118 (
            .O(N__37243),
            .I(N__37237));
    Span4Mux_v I__9117 (
            .O(N__37240),
            .I(N__37234));
    InMux I__9116 (
            .O(N__37237),
            .I(N__37231));
    Odrv4 I__9115 (
            .O(N__37234),
            .I(M_this_ext_address_qZ0Z_10));
    LocalMux I__9114 (
            .O(N__37231),
            .I(M_this_ext_address_qZ0Z_10));
    InMux I__9113 (
            .O(N__37226),
            .I(un1_M_this_ext_address_q_cry_9));
    IoInMux I__9112 (
            .O(N__37223),
            .I(N__37220));
    LocalMux I__9111 (
            .O(N__37220),
            .I(N__37217));
    IoSpan4Mux I__9110 (
            .O(N__37217),
            .I(N__37214));
    IoSpan4Mux I__9109 (
            .O(N__37214),
            .I(N__37211));
    Span4Mux_s3_v I__9108 (
            .O(N__37211),
            .I(N__37207));
    CascadeMux I__9107 (
            .O(N__37210),
            .I(N__37204));
    Span4Mux_v I__9106 (
            .O(N__37207),
            .I(N__37201));
    InMux I__9105 (
            .O(N__37204),
            .I(N__37198));
    Odrv4 I__9104 (
            .O(N__37201),
            .I(M_this_ext_address_qZ0Z_11));
    LocalMux I__9103 (
            .O(N__37198),
            .I(M_this_ext_address_qZ0Z_11));
    InMux I__9102 (
            .O(N__37193),
            .I(un1_M_this_ext_address_q_cry_10));
    IoInMux I__9101 (
            .O(N__37190),
            .I(N__37187));
    LocalMux I__9100 (
            .O(N__37187),
            .I(N__37184));
    Span4Mux_s3_h I__9099 (
            .O(N__37184),
            .I(N__37181));
    Span4Mux_h I__9098 (
            .O(N__37181),
            .I(N__37177));
    CascadeMux I__9097 (
            .O(N__37180),
            .I(N__37174));
    Span4Mux_h I__9096 (
            .O(N__37177),
            .I(N__37171));
    InMux I__9095 (
            .O(N__37174),
            .I(N__37168));
    Odrv4 I__9094 (
            .O(N__37171),
            .I(M_this_ext_address_qZ0Z_12));
    LocalMux I__9093 (
            .O(N__37168),
            .I(M_this_ext_address_qZ0Z_12));
    InMux I__9092 (
            .O(N__37163),
            .I(un1_M_this_ext_address_q_cry_11));
    IoInMux I__9091 (
            .O(N__37160),
            .I(N__37157));
    LocalMux I__9090 (
            .O(N__37157),
            .I(N__37154));
    Span4Mux_s2_h I__9089 (
            .O(N__37154),
            .I(N__37151));
    Span4Mux_v I__9088 (
            .O(N__37151),
            .I(N__37147));
    CascadeMux I__9087 (
            .O(N__37150),
            .I(N__37144));
    Sp12to4 I__9086 (
            .O(N__37147),
            .I(N__37141));
    InMux I__9085 (
            .O(N__37144),
            .I(N__37138));
    Odrv12 I__9084 (
            .O(N__37141),
            .I(M_this_ext_address_qZ0Z_13));
    LocalMux I__9083 (
            .O(N__37138),
            .I(M_this_ext_address_qZ0Z_13));
    InMux I__9082 (
            .O(N__37133),
            .I(un1_M_this_ext_address_q_cry_12));
    IoInMux I__9081 (
            .O(N__37130),
            .I(N__37127));
    LocalMux I__9080 (
            .O(N__37127),
            .I(N__37124));
    IoSpan4Mux I__9079 (
            .O(N__37124),
            .I(N__37121));
    Span4Mux_s2_h I__9078 (
            .O(N__37121),
            .I(N__37118));
    Sp12to4 I__9077 (
            .O(N__37118),
            .I(N__37114));
    CascadeMux I__9076 (
            .O(N__37117),
            .I(N__37111));
    Span12Mux_s11_h I__9075 (
            .O(N__37114),
            .I(N__37108));
    InMux I__9074 (
            .O(N__37111),
            .I(N__37105));
    Odrv12 I__9073 (
            .O(N__37108),
            .I(M_this_ext_address_qZ0Z_14));
    LocalMux I__9072 (
            .O(N__37105),
            .I(M_this_ext_address_qZ0Z_14));
    InMux I__9071 (
            .O(N__37100),
            .I(un1_M_this_ext_address_q_cry_13));
    InMux I__9070 (
            .O(N__37097),
            .I(N__37073));
    InMux I__9069 (
            .O(N__37096),
            .I(N__37073));
    InMux I__9068 (
            .O(N__37095),
            .I(N__37073));
    InMux I__9067 (
            .O(N__37094),
            .I(N__37073));
    InMux I__9066 (
            .O(N__37093),
            .I(N__37064));
    InMux I__9065 (
            .O(N__37092),
            .I(N__37064));
    InMux I__9064 (
            .O(N__37091),
            .I(N__37064));
    InMux I__9063 (
            .O(N__37090),
            .I(N__37064));
    InMux I__9062 (
            .O(N__37089),
            .I(N__37055));
    InMux I__9061 (
            .O(N__37088),
            .I(N__37055));
    InMux I__9060 (
            .O(N__37087),
            .I(N__37055));
    InMux I__9059 (
            .O(N__37086),
            .I(N__37055));
    InMux I__9058 (
            .O(N__37085),
            .I(N__37046));
    InMux I__9057 (
            .O(N__37084),
            .I(N__37046));
    InMux I__9056 (
            .O(N__37083),
            .I(N__37046));
    InMux I__9055 (
            .O(N__37082),
            .I(N__37046));
    LocalMux I__9054 (
            .O(N__37073),
            .I(N__37036));
    LocalMux I__9053 (
            .O(N__37064),
            .I(N__37036));
    LocalMux I__9052 (
            .O(N__37055),
            .I(N__37036));
    LocalMux I__9051 (
            .O(N__37046),
            .I(N__37036));
    InMux I__9050 (
            .O(N__37045),
            .I(N__37033));
    Span4Mux_v I__9049 (
            .O(N__37036),
            .I(N__37028));
    LocalMux I__9048 (
            .O(N__37033),
            .I(N__37028));
    Span4Mux_h I__9047 (
            .O(N__37028),
            .I(N__37025));
    Odrv4 I__9046 (
            .O(N__37025),
            .I(N_295));
    InMux I__9045 (
            .O(N__37022),
            .I(un1_M_this_ext_address_q_cry_14));
    IoInMux I__9044 (
            .O(N__37019),
            .I(N__37016));
    LocalMux I__9043 (
            .O(N__37016),
            .I(N__37013));
    Span4Mux_s2_h I__9042 (
            .O(N__37013),
            .I(N__37010));
    Sp12to4 I__9041 (
            .O(N__37010),
            .I(N__37007));
    Span12Mux_v I__9040 (
            .O(N__37007),
            .I(N__37004));
    Span12Mux_v I__9039 (
            .O(N__37004),
            .I(N__37000));
    InMux I__9038 (
            .O(N__37003),
            .I(N__36997));
    Odrv12 I__9037 (
            .O(N__37000),
            .I(M_this_ext_address_qZ0Z_15));
    LocalMux I__9036 (
            .O(N__36997),
            .I(M_this_ext_address_qZ0Z_15));
    CascadeMux I__9035 (
            .O(N__36992),
            .I(N__36988));
    CascadeMux I__9034 (
            .O(N__36991),
            .I(N__36985));
    InMux I__9033 (
            .O(N__36988),
            .I(N__36979));
    InMux I__9032 (
            .O(N__36985),
            .I(N__36979));
    CascadeMux I__9031 (
            .O(N__36984),
            .I(N__36976));
    LocalMux I__9030 (
            .O(N__36979),
            .I(N__36973));
    InMux I__9029 (
            .O(N__36976),
            .I(N__36970));
    Odrv4 I__9028 (
            .O(N__36973),
            .I(\this_start_data_delay.N_231_0 ));
    LocalMux I__9027 (
            .O(N__36970),
            .I(\this_start_data_delay.N_231_0 ));
    CascadeMux I__9026 (
            .O(N__36965),
            .I(N__36944));
    CascadeMux I__9025 (
            .O(N__36964),
            .I(N__36940));
    CascadeMux I__9024 (
            .O(N__36963),
            .I(N__36930));
    InMux I__9023 (
            .O(N__36962),
            .I(N__36922));
    InMux I__9022 (
            .O(N__36961),
            .I(N__36922));
    InMux I__9021 (
            .O(N__36960),
            .I(N__36917));
    InMux I__9020 (
            .O(N__36959),
            .I(N__36917));
    InMux I__9019 (
            .O(N__36958),
            .I(N__36914));
    InMux I__9018 (
            .O(N__36957),
            .I(N__36911));
    InMux I__9017 (
            .O(N__36956),
            .I(N__36906));
    InMux I__9016 (
            .O(N__36955),
            .I(N__36906));
    InMux I__9015 (
            .O(N__36954),
            .I(N__36903));
    InMux I__9014 (
            .O(N__36953),
            .I(N__36898));
    InMux I__9013 (
            .O(N__36952),
            .I(N__36898));
    InMux I__9012 (
            .O(N__36951),
            .I(N__36895));
    InMux I__9011 (
            .O(N__36950),
            .I(N__36892));
    InMux I__9010 (
            .O(N__36949),
            .I(N__36887));
    InMux I__9009 (
            .O(N__36948),
            .I(N__36887));
    InMux I__9008 (
            .O(N__36947),
            .I(N__36884));
    InMux I__9007 (
            .O(N__36944),
            .I(N__36881));
    InMux I__9006 (
            .O(N__36943),
            .I(N__36878));
    InMux I__9005 (
            .O(N__36940),
            .I(N__36875));
    InMux I__9004 (
            .O(N__36939),
            .I(N__36868));
    InMux I__9003 (
            .O(N__36938),
            .I(N__36868));
    InMux I__9002 (
            .O(N__36937),
            .I(N__36868));
    InMux I__9001 (
            .O(N__36936),
            .I(N__36865));
    InMux I__9000 (
            .O(N__36935),
            .I(N__36862));
    InMux I__8999 (
            .O(N__36934),
            .I(N__36859));
    InMux I__8998 (
            .O(N__36933),
            .I(N__36856));
    InMux I__8997 (
            .O(N__36930),
            .I(N__36851));
    InMux I__8996 (
            .O(N__36929),
            .I(N__36851));
    InMux I__8995 (
            .O(N__36928),
            .I(N__36846));
    InMux I__8994 (
            .O(N__36927),
            .I(N__36846));
    LocalMux I__8993 (
            .O(N__36922),
            .I(N__36809));
    LocalMux I__8992 (
            .O(N__36917),
            .I(N__36806));
    LocalMux I__8991 (
            .O(N__36914),
            .I(N__36803));
    LocalMux I__8990 (
            .O(N__36911),
            .I(N__36800));
    LocalMux I__8989 (
            .O(N__36906),
            .I(N__36797));
    LocalMux I__8988 (
            .O(N__36903),
            .I(N__36794));
    LocalMux I__8987 (
            .O(N__36898),
            .I(N__36791));
    LocalMux I__8986 (
            .O(N__36895),
            .I(N__36788));
    LocalMux I__8985 (
            .O(N__36892),
            .I(N__36785));
    LocalMux I__8984 (
            .O(N__36887),
            .I(N__36782));
    LocalMux I__8983 (
            .O(N__36884),
            .I(N__36779));
    LocalMux I__8982 (
            .O(N__36881),
            .I(N__36776));
    LocalMux I__8981 (
            .O(N__36878),
            .I(N__36773));
    LocalMux I__8980 (
            .O(N__36875),
            .I(N__36770));
    LocalMux I__8979 (
            .O(N__36868),
            .I(N__36767));
    LocalMux I__8978 (
            .O(N__36865),
            .I(N__36764));
    LocalMux I__8977 (
            .O(N__36862),
            .I(N__36761));
    LocalMux I__8976 (
            .O(N__36859),
            .I(N__36758));
    LocalMux I__8975 (
            .O(N__36856),
            .I(N__36755));
    LocalMux I__8974 (
            .O(N__36851),
            .I(N__36752));
    LocalMux I__8973 (
            .O(N__36846),
            .I(N__36749));
    SRMux I__8972 (
            .O(N__36845),
            .I(N__36638));
    SRMux I__8971 (
            .O(N__36844),
            .I(N__36638));
    SRMux I__8970 (
            .O(N__36843),
            .I(N__36638));
    SRMux I__8969 (
            .O(N__36842),
            .I(N__36638));
    SRMux I__8968 (
            .O(N__36841),
            .I(N__36638));
    SRMux I__8967 (
            .O(N__36840),
            .I(N__36638));
    SRMux I__8966 (
            .O(N__36839),
            .I(N__36638));
    SRMux I__8965 (
            .O(N__36838),
            .I(N__36638));
    SRMux I__8964 (
            .O(N__36837),
            .I(N__36638));
    SRMux I__8963 (
            .O(N__36836),
            .I(N__36638));
    SRMux I__8962 (
            .O(N__36835),
            .I(N__36638));
    SRMux I__8961 (
            .O(N__36834),
            .I(N__36638));
    SRMux I__8960 (
            .O(N__36833),
            .I(N__36638));
    SRMux I__8959 (
            .O(N__36832),
            .I(N__36638));
    SRMux I__8958 (
            .O(N__36831),
            .I(N__36638));
    SRMux I__8957 (
            .O(N__36830),
            .I(N__36638));
    SRMux I__8956 (
            .O(N__36829),
            .I(N__36638));
    SRMux I__8955 (
            .O(N__36828),
            .I(N__36638));
    SRMux I__8954 (
            .O(N__36827),
            .I(N__36638));
    SRMux I__8953 (
            .O(N__36826),
            .I(N__36638));
    SRMux I__8952 (
            .O(N__36825),
            .I(N__36638));
    SRMux I__8951 (
            .O(N__36824),
            .I(N__36638));
    SRMux I__8950 (
            .O(N__36823),
            .I(N__36638));
    SRMux I__8949 (
            .O(N__36822),
            .I(N__36638));
    SRMux I__8948 (
            .O(N__36821),
            .I(N__36638));
    SRMux I__8947 (
            .O(N__36820),
            .I(N__36638));
    SRMux I__8946 (
            .O(N__36819),
            .I(N__36638));
    SRMux I__8945 (
            .O(N__36818),
            .I(N__36638));
    SRMux I__8944 (
            .O(N__36817),
            .I(N__36638));
    SRMux I__8943 (
            .O(N__36816),
            .I(N__36638));
    SRMux I__8942 (
            .O(N__36815),
            .I(N__36638));
    SRMux I__8941 (
            .O(N__36814),
            .I(N__36638));
    SRMux I__8940 (
            .O(N__36813),
            .I(N__36638));
    SRMux I__8939 (
            .O(N__36812),
            .I(N__36638));
    Glb2LocalMux I__8938 (
            .O(N__36809),
            .I(N__36638));
    Glb2LocalMux I__8937 (
            .O(N__36806),
            .I(N__36638));
    Glb2LocalMux I__8936 (
            .O(N__36803),
            .I(N__36638));
    Glb2LocalMux I__8935 (
            .O(N__36800),
            .I(N__36638));
    Glb2LocalMux I__8934 (
            .O(N__36797),
            .I(N__36638));
    Glb2LocalMux I__8933 (
            .O(N__36794),
            .I(N__36638));
    Glb2LocalMux I__8932 (
            .O(N__36791),
            .I(N__36638));
    Glb2LocalMux I__8931 (
            .O(N__36788),
            .I(N__36638));
    Glb2LocalMux I__8930 (
            .O(N__36785),
            .I(N__36638));
    Glb2LocalMux I__8929 (
            .O(N__36782),
            .I(N__36638));
    Glb2LocalMux I__8928 (
            .O(N__36779),
            .I(N__36638));
    Glb2LocalMux I__8927 (
            .O(N__36776),
            .I(N__36638));
    Glb2LocalMux I__8926 (
            .O(N__36773),
            .I(N__36638));
    Glb2LocalMux I__8925 (
            .O(N__36770),
            .I(N__36638));
    Glb2LocalMux I__8924 (
            .O(N__36767),
            .I(N__36638));
    Glb2LocalMux I__8923 (
            .O(N__36764),
            .I(N__36638));
    Glb2LocalMux I__8922 (
            .O(N__36761),
            .I(N__36638));
    Glb2LocalMux I__8921 (
            .O(N__36758),
            .I(N__36638));
    Glb2LocalMux I__8920 (
            .O(N__36755),
            .I(N__36638));
    Glb2LocalMux I__8919 (
            .O(N__36752),
            .I(N__36638));
    Glb2LocalMux I__8918 (
            .O(N__36749),
            .I(N__36638));
    GlobalMux I__8917 (
            .O(N__36638),
            .I(N__36635));
    gio2CtrlBuf I__8916 (
            .O(N__36635),
            .I(M_this_reset_cond_out_g_0));
    InMux I__8915 (
            .O(N__36632),
            .I(N__36626));
    InMux I__8914 (
            .O(N__36631),
            .I(N__36623));
    InMux I__8913 (
            .O(N__36630),
            .I(N__36618));
    InMux I__8912 (
            .O(N__36629),
            .I(N__36618));
    LocalMux I__8911 (
            .O(N__36626),
            .I(N__36609));
    LocalMux I__8910 (
            .O(N__36623),
            .I(N__36609));
    LocalMux I__8909 (
            .O(N__36618),
            .I(N__36609));
    InMux I__8908 (
            .O(N__36617),
            .I(N__36604));
    InMux I__8907 (
            .O(N__36616),
            .I(N__36604));
    Span12Mux_h I__8906 (
            .O(N__36609),
            .I(N__36599));
    LocalMux I__8905 (
            .O(N__36604),
            .I(N__36599));
    Span12Mux_v I__8904 (
            .O(N__36599),
            .I(N__36596));
    Odrv12 I__8903 (
            .O(N__36596),
            .I(\this_start_data_delay.N_227_0 ));
    InMux I__8902 (
            .O(N__36593),
            .I(N__36588));
    InMux I__8901 (
            .O(N__36592),
            .I(N__36583));
    InMux I__8900 (
            .O(N__36591),
            .I(N__36583));
    LocalMux I__8899 (
            .O(N__36588),
            .I(N__36580));
    LocalMux I__8898 (
            .O(N__36583),
            .I(\this_start_data_delay.N_242_0 ));
    Odrv4 I__8897 (
            .O(N__36580),
            .I(\this_start_data_delay.N_242_0 ));
    CascadeMux I__8896 (
            .O(N__36575),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_ ));
    CascadeMux I__8895 (
            .O(N__36572),
            .I(N__36569));
    InMux I__8894 (
            .O(N__36569),
            .I(N__36559));
    InMux I__8893 (
            .O(N__36568),
            .I(N__36556));
    InMux I__8892 (
            .O(N__36567),
            .I(N__36553));
    CascadeMux I__8891 (
            .O(N__36566),
            .I(N__36547));
    InMux I__8890 (
            .O(N__36565),
            .I(N__36540));
    InMux I__8889 (
            .O(N__36564),
            .I(N__36532));
    InMux I__8888 (
            .O(N__36563),
            .I(N__36532));
    InMux I__8887 (
            .O(N__36562),
            .I(N__36532));
    LocalMux I__8886 (
            .O(N__36559),
            .I(N__36527));
    LocalMux I__8885 (
            .O(N__36556),
            .I(N__36527));
    LocalMux I__8884 (
            .O(N__36553),
            .I(N__36524));
    InMux I__8883 (
            .O(N__36552),
            .I(N__36521));
    InMux I__8882 (
            .O(N__36551),
            .I(N__36518));
    InMux I__8881 (
            .O(N__36550),
            .I(N__36515));
    InMux I__8880 (
            .O(N__36547),
            .I(N__36512));
    InMux I__8879 (
            .O(N__36546),
            .I(N__36509));
    InMux I__8878 (
            .O(N__36545),
            .I(N__36506));
    InMux I__8877 (
            .O(N__36544),
            .I(N__36503));
    InMux I__8876 (
            .O(N__36543),
            .I(N__36499));
    LocalMux I__8875 (
            .O(N__36540),
            .I(N__36495));
    InMux I__8874 (
            .O(N__36539),
            .I(N__36491));
    LocalMux I__8873 (
            .O(N__36532),
            .I(N__36486));
    Span4Mux_v I__8872 (
            .O(N__36527),
            .I(N__36486));
    Span4Mux_v I__8871 (
            .O(N__36524),
            .I(N__36483));
    LocalMux I__8870 (
            .O(N__36521),
            .I(N__36474));
    LocalMux I__8869 (
            .O(N__36518),
            .I(N__36474));
    LocalMux I__8868 (
            .O(N__36515),
            .I(N__36474));
    LocalMux I__8867 (
            .O(N__36512),
            .I(N__36474));
    LocalMux I__8866 (
            .O(N__36509),
            .I(N__36469));
    LocalMux I__8865 (
            .O(N__36506),
            .I(N__36469));
    LocalMux I__8864 (
            .O(N__36503),
            .I(N__36466));
    InMux I__8863 (
            .O(N__36502),
            .I(N__36463));
    LocalMux I__8862 (
            .O(N__36499),
            .I(N__36460));
    InMux I__8861 (
            .O(N__36498),
            .I(N__36457));
    Span4Mux_h I__8860 (
            .O(N__36495),
            .I(N__36454));
    InMux I__8859 (
            .O(N__36494),
            .I(N__36451));
    LocalMux I__8858 (
            .O(N__36491),
            .I(N__36448));
    Span4Mux_h I__8857 (
            .O(N__36486),
            .I(N__36439));
    Span4Mux_v I__8856 (
            .O(N__36483),
            .I(N__36439));
    Span4Mux_v I__8855 (
            .O(N__36474),
            .I(N__36439));
    Span4Mux_v I__8854 (
            .O(N__36469),
            .I(N__36439));
    Odrv4 I__8853 (
            .O(N__36466),
            .I(N_220_0));
    LocalMux I__8852 (
            .O(N__36463),
            .I(N_220_0));
    Odrv12 I__8851 (
            .O(N__36460),
            .I(N_220_0));
    LocalMux I__8850 (
            .O(N__36457),
            .I(N_220_0));
    Odrv4 I__8849 (
            .O(N__36454),
            .I(N_220_0));
    LocalMux I__8848 (
            .O(N__36451),
            .I(N_220_0));
    Odrv12 I__8847 (
            .O(N__36448),
            .I(N_220_0));
    Odrv4 I__8846 (
            .O(N__36439),
            .I(N_220_0));
    CascadeMux I__8845 (
            .O(N__36422),
            .I(N__36418));
    InMux I__8844 (
            .O(N__36421),
            .I(N__36415));
    InMux I__8843 (
            .O(N__36418),
            .I(N__36410));
    LocalMux I__8842 (
            .O(N__36415),
            .I(N__36407));
    InMux I__8841 (
            .O(N__36414),
            .I(N__36404));
    InMux I__8840 (
            .O(N__36413),
            .I(N__36401));
    LocalMux I__8839 (
            .O(N__36410),
            .I(M_this_state_qZ0Z_10));
    Odrv4 I__8838 (
            .O(N__36407),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__8837 (
            .O(N__36404),
            .I(M_this_state_qZ0Z_10));
    LocalMux I__8836 (
            .O(N__36401),
            .I(M_this_state_qZ0Z_10));
    IoInMux I__8835 (
            .O(N__36392),
            .I(N__36389));
    LocalMux I__8834 (
            .O(N__36389),
            .I(N__36386));
    Span4Mux_s1_v I__8833 (
            .O(N__36386),
            .I(N__36383));
    Span4Mux_v I__8832 (
            .O(N__36383),
            .I(N__36379));
    InMux I__8831 (
            .O(N__36382),
            .I(N__36376));
    Odrv4 I__8830 (
            .O(N__36379),
            .I(M_this_ext_address_qZ0Z_2));
    LocalMux I__8829 (
            .O(N__36376),
            .I(M_this_ext_address_qZ0Z_2));
    InMux I__8828 (
            .O(N__36371),
            .I(un1_M_this_ext_address_q_cry_1));
    IoInMux I__8827 (
            .O(N__36368),
            .I(N__36365));
    LocalMux I__8826 (
            .O(N__36365),
            .I(N__36362));
    Span4Mux_s3_h I__8825 (
            .O(N__36362),
            .I(N__36359));
    Span4Mux_h I__8824 (
            .O(N__36359),
            .I(N__36356));
    Span4Mux_v I__8823 (
            .O(N__36356),
            .I(N__36352));
    InMux I__8822 (
            .O(N__36355),
            .I(N__36349));
    Odrv4 I__8821 (
            .O(N__36352),
            .I(M_this_ext_address_qZ0Z_3));
    LocalMux I__8820 (
            .O(N__36349),
            .I(M_this_ext_address_qZ0Z_3));
    InMux I__8819 (
            .O(N__36344),
            .I(un1_M_this_ext_address_q_cry_2));
    IoInMux I__8818 (
            .O(N__36341),
            .I(N__36338));
    LocalMux I__8817 (
            .O(N__36338),
            .I(N__36335));
    Span4Mux_s3_h I__8816 (
            .O(N__36335),
            .I(N__36332));
    Span4Mux_h I__8815 (
            .O(N__36332),
            .I(N__36329));
    Span4Mux_h I__8814 (
            .O(N__36329),
            .I(N__36325));
    InMux I__8813 (
            .O(N__36328),
            .I(N__36322));
    Odrv4 I__8812 (
            .O(N__36325),
            .I(M_this_ext_address_qZ0Z_4));
    LocalMux I__8811 (
            .O(N__36322),
            .I(M_this_ext_address_qZ0Z_4));
    InMux I__8810 (
            .O(N__36317),
            .I(un1_M_this_ext_address_q_cry_3));
    IoInMux I__8809 (
            .O(N__36314),
            .I(N__36311));
    LocalMux I__8808 (
            .O(N__36311),
            .I(N__36308));
    IoSpan4Mux I__8807 (
            .O(N__36308),
            .I(N__36305));
    Span4Mux_s3_h I__8806 (
            .O(N__36305),
            .I(N__36302));
    Span4Mux_h I__8805 (
            .O(N__36302),
            .I(N__36298));
    InMux I__8804 (
            .O(N__36301),
            .I(N__36295));
    Odrv4 I__8803 (
            .O(N__36298),
            .I(M_this_ext_address_qZ0Z_5));
    LocalMux I__8802 (
            .O(N__36295),
            .I(M_this_ext_address_qZ0Z_5));
    InMux I__8801 (
            .O(N__36290),
            .I(un1_M_this_ext_address_q_cry_4));
    IoInMux I__8800 (
            .O(N__36287),
            .I(N__36284));
    LocalMux I__8799 (
            .O(N__36284),
            .I(N__36281));
    IoSpan4Mux I__8798 (
            .O(N__36281),
            .I(N__36278));
    IoSpan4Mux I__8797 (
            .O(N__36278),
            .I(N__36275));
    Span4Mux_s0_h I__8796 (
            .O(N__36275),
            .I(N__36272));
    Sp12to4 I__8795 (
            .O(N__36272),
            .I(N__36268));
    InMux I__8794 (
            .O(N__36271),
            .I(N__36265));
    Odrv12 I__8793 (
            .O(N__36268),
            .I(M_this_ext_address_qZ0Z_6));
    LocalMux I__8792 (
            .O(N__36265),
            .I(M_this_ext_address_qZ0Z_6));
    InMux I__8791 (
            .O(N__36260),
            .I(un1_M_this_ext_address_q_cry_5));
    IoInMux I__8790 (
            .O(N__36257),
            .I(N__36254));
    LocalMux I__8789 (
            .O(N__36254),
            .I(N__36251));
    Span4Mux_s2_h I__8788 (
            .O(N__36251),
            .I(N__36248));
    Sp12to4 I__8787 (
            .O(N__36248),
            .I(N__36245));
    Span12Mux_s11_v I__8786 (
            .O(N__36245),
            .I(N__36242));
    Span12Mux_v I__8785 (
            .O(N__36242),
            .I(N__36238));
    InMux I__8784 (
            .O(N__36241),
            .I(N__36235));
    Odrv12 I__8783 (
            .O(N__36238),
            .I(M_this_ext_address_qZ0Z_7));
    LocalMux I__8782 (
            .O(N__36235),
            .I(M_this_ext_address_qZ0Z_7));
    InMux I__8781 (
            .O(N__36230),
            .I(un1_M_this_ext_address_q_cry_6));
    IoInMux I__8780 (
            .O(N__36227),
            .I(N__36224));
    LocalMux I__8779 (
            .O(N__36224),
            .I(N__36221));
    IoSpan4Mux I__8778 (
            .O(N__36221),
            .I(N__36218));
    Span4Mux_s3_v I__8777 (
            .O(N__36218),
            .I(N__36214));
    CascadeMux I__8776 (
            .O(N__36217),
            .I(N__36211));
    Span4Mux_v I__8775 (
            .O(N__36214),
            .I(N__36208));
    InMux I__8774 (
            .O(N__36211),
            .I(N__36205));
    Odrv4 I__8773 (
            .O(N__36208),
            .I(M_this_ext_address_qZ0Z_8));
    LocalMux I__8772 (
            .O(N__36205),
            .I(M_this_ext_address_qZ0Z_8));
    InMux I__8771 (
            .O(N__36200),
            .I(bfn_21_25_0_));
    IoInMux I__8770 (
            .O(N__36197),
            .I(N__36194));
    LocalMux I__8769 (
            .O(N__36194),
            .I(N__36191));
    Span4Mux_s3_v I__8768 (
            .O(N__36191),
            .I(N__36187));
    CascadeMux I__8767 (
            .O(N__36190),
            .I(N__36184));
    Span4Mux_v I__8766 (
            .O(N__36187),
            .I(N__36181));
    InMux I__8765 (
            .O(N__36184),
            .I(N__36178));
    Odrv4 I__8764 (
            .O(N__36181),
            .I(M_this_ext_address_qZ0Z_9));
    LocalMux I__8763 (
            .O(N__36178),
            .I(M_this_ext_address_qZ0Z_9));
    InMux I__8762 (
            .O(N__36173),
            .I(un1_M_this_ext_address_q_cry_8));
    InMux I__8761 (
            .O(N__36170),
            .I(N__36167));
    LocalMux I__8760 (
            .O(N__36167),
            .I(N__36162));
    InMux I__8759 (
            .O(N__36166),
            .I(N__36157));
    InMux I__8758 (
            .O(N__36165),
            .I(N__36154));
    Span12Mux_h I__8757 (
            .O(N__36162),
            .I(N__36151));
    InMux I__8756 (
            .O(N__36161),
            .I(N__36148));
    InMux I__8755 (
            .O(N__36160),
            .I(N__36145));
    LocalMux I__8754 (
            .O(N__36157),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__8753 (
            .O(N__36154),
            .I(M_this_state_qZ0Z_6));
    Odrv12 I__8752 (
            .O(N__36151),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__8751 (
            .O(N__36148),
            .I(M_this_state_qZ0Z_6));
    LocalMux I__8750 (
            .O(N__36145),
            .I(M_this_state_qZ0Z_6));
    InMux I__8749 (
            .O(N__36134),
            .I(N__36131));
    LocalMux I__8748 (
            .O(N__36131),
            .I(N__36127));
    InMux I__8747 (
            .O(N__36130),
            .I(N__36122));
    Span4Mux_h I__8746 (
            .O(N__36127),
            .I(N__36119));
    InMux I__8745 (
            .O(N__36126),
            .I(N__36114));
    InMux I__8744 (
            .O(N__36125),
            .I(N__36114));
    LocalMux I__8743 (
            .O(N__36122),
            .I(N__36111));
    Odrv4 I__8742 (
            .O(N__36119),
            .I(M_this_state_qZ0Z_5));
    LocalMux I__8741 (
            .O(N__36114),
            .I(M_this_state_qZ0Z_5));
    Odrv4 I__8740 (
            .O(N__36111),
            .I(M_this_state_qZ0Z_5));
    InMux I__8739 (
            .O(N__36104),
            .I(N__36101));
    LocalMux I__8738 (
            .O(N__36101),
            .I(N__36098));
    Span4Mux_h I__8737 (
            .O(N__36098),
            .I(N__36094));
    InMux I__8736 (
            .O(N__36097),
            .I(N__36091));
    Odrv4 I__8735 (
            .O(N__36094),
            .I(\this_start_data_delay.N_239_0 ));
    LocalMux I__8734 (
            .O(N__36091),
            .I(\this_start_data_delay.N_239_0 ));
    InMux I__8733 (
            .O(N__36086),
            .I(N__36080));
    InMux I__8732 (
            .O(N__36085),
            .I(N__36077));
    InMux I__8731 (
            .O(N__36084),
            .I(N__36072));
    InMux I__8730 (
            .O(N__36083),
            .I(N__36072));
    LocalMux I__8729 (
            .O(N__36080),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__8728 (
            .O(N__36077),
            .I(M_this_state_qZ0Z_3));
    LocalMux I__8727 (
            .O(N__36072),
            .I(M_this_state_qZ0Z_3));
    InMux I__8726 (
            .O(N__36065),
            .I(N__36062));
    LocalMux I__8725 (
            .O(N__36062),
            .I(N__36059));
    Span4Mux_h I__8724 (
            .O(N__36059),
            .I(N__36056));
    Span4Mux_h I__8723 (
            .O(N__36056),
            .I(N__36050));
    InMux I__8722 (
            .O(N__36055),
            .I(N__36047));
    InMux I__8721 (
            .O(N__36054),
            .I(N__36042));
    InMux I__8720 (
            .O(N__36053),
            .I(N__36042));
    Odrv4 I__8719 (
            .O(N__36050),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__8718 (
            .O(N__36047),
            .I(M_this_state_qZ0Z_2));
    LocalMux I__8717 (
            .O(N__36042),
            .I(M_this_state_qZ0Z_2));
    CascadeMux I__8716 (
            .O(N__36035),
            .I(N__36029));
    InMux I__8715 (
            .O(N__36034),
            .I(N__36024));
    InMux I__8714 (
            .O(N__36033),
            .I(N__36024));
    InMux I__8713 (
            .O(N__36032),
            .I(N__36021));
    InMux I__8712 (
            .O(N__36029),
            .I(N__36017));
    LocalMux I__8711 (
            .O(N__36024),
            .I(N__36014));
    LocalMux I__8710 (
            .O(N__36021),
            .I(N__36011));
    InMux I__8709 (
            .O(N__36020),
            .I(N__36008));
    LocalMux I__8708 (
            .O(N__36017),
            .I(N__36002));
    Span4Mux_v I__8707 (
            .O(N__36014),
            .I(N__36002));
    Span12Mux_v I__8706 (
            .O(N__36011),
            .I(N__35999));
    LocalMux I__8705 (
            .O(N__36008),
            .I(N__35996));
    InMux I__8704 (
            .O(N__36007),
            .I(N__35993));
    Odrv4 I__8703 (
            .O(N__36002),
            .I(M_this_state_qZ0Z_1));
    Odrv12 I__8702 (
            .O(N__35999),
            .I(M_this_state_qZ0Z_1));
    Odrv4 I__8701 (
            .O(N__35996),
            .I(M_this_state_qZ0Z_1));
    LocalMux I__8700 (
            .O(N__35993),
            .I(M_this_state_qZ0Z_1));
    InMux I__8699 (
            .O(N__35984),
            .I(N__35980));
    InMux I__8698 (
            .O(N__35983),
            .I(N__35977));
    LocalMux I__8697 (
            .O(N__35980),
            .I(\this_start_data_delay.N_420_3 ));
    LocalMux I__8696 (
            .O(N__35977),
            .I(\this_start_data_delay.N_420_3 ));
    InMux I__8695 (
            .O(N__35972),
            .I(N__35966));
    InMux I__8694 (
            .O(N__35971),
            .I(N__35966));
    LocalMux I__8693 (
            .O(N__35966),
            .I(N__35957));
    InMux I__8692 (
            .O(N__35965),
            .I(N__35954));
    InMux I__8691 (
            .O(N__35964),
            .I(N__35951));
    InMux I__8690 (
            .O(N__35963),
            .I(N__35948));
    InMux I__8689 (
            .O(N__35962),
            .I(N__35945));
    InMux I__8688 (
            .O(N__35961),
            .I(N__35942));
    InMux I__8687 (
            .O(N__35960),
            .I(N__35939));
    Odrv4 I__8686 (
            .O(N__35957),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8685 (
            .O(N__35954),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8684 (
            .O(N__35951),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8683 (
            .O(N__35948),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8682 (
            .O(N__35945),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8681 (
            .O(N__35942),
            .I(\this_start_data_delay.N_23_1_0 ));
    LocalMux I__8680 (
            .O(N__35939),
            .I(\this_start_data_delay.N_23_1_0 ));
    CascadeMux I__8679 (
            .O(N__35924),
            .I(\this_start_data_delay.N_344_cascade_ ));
    InMux I__8678 (
            .O(N__35921),
            .I(N__35917));
    InMux I__8677 (
            .O(N__35920),
            .I(N__35914));
    LocalMux I__8676 (
            .O(N__35917),
            .I(N_465));
    LocalMux I__8675 (
            .O(N__35914),
            .I(N_465));
    InMux I__8674 (
            .O(N__35909),
            .I(N__35906));
    LocalMux I__8673 (
            .O(N__35906),
            .I(N__35901));
    InMux I__8672 (
            .O(N__35905),
            .I(N__35896));
    InMux I__8671 (
            .O(N__35904),
            .I(N__35896));
    Span4Mux_h I__8670 (
            .O(N__35901),
            .I(N__35893));
    LocalMux I__8669 (
            .O(N__35896),
            .I(N__35890));
    Odrv4 I__8668 (
            .O(N__35893),
            .I(\this_start_data_delay.N_246_0 ));
    Odrv4 I__8667 (
            .O(N__35890),
            .I(\this_start_data_delay.N_246_0 ));
    InMux I__8666 (
            .O(N__35885),
            .I(N__35882));
    LocalMux I__8665 (
            .O(N__35882),
            .I(\this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0 ));
    CascadeMux I__8664 (
            .O(N__35879),
            .I(N__35875));
    InMux I__8663 (
            .O(N__35878),
            .I(N__35872));
    InMux I__8662 (
            .O(N__35875),
            .I(N__35869));
    LocalMux I__8661 (
            .O(N__35872),
            .I(N__35864));
    LocalMux I__8660 (
            .O(N__35869),
            .I(N__35864));
    Span4Mux_v I__8659 (
            .O(N__35864),
            .I(N__35861));
    Odrv4 I__8658 (
            .O(N__35861),
            .I(M_last_q_RNIE8SF1));
    IoInMux I__8657 (
            .O(N__35858),
            .I(N__35855));
    LocalMux I__8656 (
            .O(N__35855),
            .I(N__35852));
    Span12Mux_s8_v I__8655 (
            .O(N__35852),
            .I(N__35848));
    InMux I__8654 (
            .O(N__35851),
            .I(N__35845));
    Odrv12 I__8653 (
            .O(N__35848),
            .I(M_this_ext_address_qZ0Z_0));
    LocalMux I__8652 (
            .O(N__35845),
            .I(M_this_ext_address_qZ0Z_0));
    IoInMux I__8651 (
            .O(N__35840),
            .I(N__35837));
    LocalMux I__8650 (
            .O(N__35837),
            .I(N__35834));
    Span4Mux_s2_v I__8649 (
            .O(N__35834),
            .I(N__35831));
    Span4Mux_h I__8648 (
            .O(N__35831),
            .I(N__35828));
    Span4Mux_v I__8647 (
            .O(N__35828),
            .I(N__35824));
    InMux I__8646 (
            .O(N__35827),
            .I(N__35821));
    Odrv4 I__8645 (
            .O(N__35824),
            .I(M_this_ext_address_qZ0Z_1));
    LocalMux I__8644 (
            .O(N__35821),
            .I(M_this_ext_address_qZ0Z_1));
    InMux I__8643 (
            .O(N__35816),
            .I(un1_M_this_ext_address_q_cry_0));
    InMux I__8642 (
            .O(N__35813),
            .I(N__35796));
    InMux I__8641 (
            .O(N__35812),
            .I(N__35796));
    InMux I__8640 (
            .O(N__35811),
            .I(N__35796));
    InMux I__8639 (
            .O(N__35810),
            .I(N__35796));
    InMux I__8638 (
            .O(N__35809),
            .I(N__35787));
    InMux I__8637 (
            .O(N__35808),
            .I(N__35787));
    InMux I__8636 (
            .O(N__35807),
            .I(N__35787));
    InMux I__8635 (
            .O(N__35806),
            .I(N__35787));
    InMux I__8634 (
            .O(N__35805),
            .I(N__35778));
    LocalMux I__8633 (
            .O(N__35796),
            .I(N__35772));
    LocalMux I__8632 (
            .O(N__35787),
            .I(N__35772));
    InMux I__8631 (
            .O(N__35786),
            .I(N__35767));
    InMux I__8630 (
            .O(N__35785),
            .I(N__35767));
    InMux I__8629 (
            .O(N__35784),
            .I(N__35758));
    InMux I__8628 (
            .O(N__35783),
            .I(N__35758));
    InMux I__8627 (
            .O(N__35782),
            .I(N__35758));
    InMux I__8626 (
            .O(N__35781),
            .I(N__35758));
    LocalMux I__8625 (
            .O(N__35778),
            .I(N__35755));
    CascadeMux I__8624 (
            .O(N__35777),
            .I(N__35752));
    Span4Mux_h I__8623 (
            .O(N__35772),
            .I(N__35745));
    LocalMux I__8622 (
            .O(N__35767),
            .I(N__35745));
    LocalMux I__8621 (
            .O(N__35758),
            .I(N__35745));
    Span4Mux_h I__8620 (
            .O(N__35755),
            .I(N__35742));
    InMux I__8619 (
            .O(N__35752),
            .I(N__35739));
    Span4Mux_v I__8618 (
            .O(N__35745),
            .I(N__35736));
    Odrv4 I__8617 (
            .O(N__35742),
            .I(N_241_0));
    LocalMux I__8616 (
            .O(N__35739),
            .I(N_241_0));
    Odrv4 I__8615 (
            .O(N__35736),
            .I(N_241_0));
    CascadeMux I__8614 (
            .O(N__35729),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_ ));
    InMux I__8613 (
            .O(N__35726),
            .I(N__35723));
    LocalMux I__8612 (
            .O(N__35723),
            .I(N__35720));
    Span4Mux_h I__8611 (
            .O(N__35720),
            .I(N__35717));
    Odrv4 I__8610 (
            .O(N__35717),
            .I(\this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0 ));
    InMux I__8609 (
            .O(N__35714),
            .I(N__35707));
    CascadeMux I__8608 (
            .O(N__35713),
            .I(N__35704));
    InMux I__8607 (
            .O(N__35712),
            .I(N__35701));
    InMux I__8606 (
            .O(N__35711),
            .I(N__35696));
    InMux I__8605 (
            .O(N__35710),
            .I(N__35696));
    LocalMux I__8604 (
            .O(N__35707),
            .I(N__35692));
    InMux I__8603 (
            .O(N__35704),
            .I(N__35689));
    LocalMux I__8602 (
            .O(N__35701),
            .I(N__35686));
    LocalMux I__8601 (
            .O(N__35696),
            .I(N__35683));
    InMux I__8600 (
            .O(N__35695),
            .I(N__35680));
    Odrv4 I__8599 (
            .O(N__35692),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__8598 (
            .O(N__35689),
            .I(M_this_state_qZ0Z_12));
    Odrv12 I__8597 (
            .O(N__35686),
            .I(M_this_state_qZ0Z_12));
    Odrv4 I__8596 (
            .O(N__35683),
            .I(M_this_state_qZ0Z_12));
    LocalMux I__8595 (
            .O(N__35680),
            .I(M_this_state_qZ0Z_12));
    CascadeMux I__8594 (
            .O(N__35669),
            .I(N__35666));
    InMux I__8593 (
            .O(N__35666),
            .I(N__35663));
    LocalMux I__8592 (
            .O(N__35663),
            .I(\this_start_data_delay.N_245_0 ));
    InMux I__8591 (
            .O(N__35660),
            .I(N__35657));
    LocalMux I__8590 (
            .O(N__35657),
            .I(N__35649));
    InMux I__8589 (
            .O(N__35656),
            .I(N__35638));
    InMux I__8588 (
            .O(N__35655),
            .I(N__35638));
    InMux I__8587 (
            .O(N__35654),
            .I(N__35638));
    InMux I__8586 (
            .O(N__35653),
            .I(N__35638));
    InMux I__8585 (
            .O(N__35652),
            .I(N__35638));
    Odrv12 I__8584 (
            .O(N__35649),
            .I(M_this_state_qZ0Z_7));
    LocalMux I__8583 (
            .O(N__35638),
            .I(M_this_state_qZ0Z_7));
    InMux I__8582 (
            .O(N__35633),
            .I(N__35630));
    LocalMux I__8581 (
            .O(N__35630),
            .I(N__35625));
    InMux I__8580 (
            .O(N__35629),
            .I(N__35622));
    InMux I__8579 (
            .O(N__35628),
            .I(N__35617));
    Span4Mux_h I__8578 (
            .O(N__35625),
            .I(N__35612));
    LocalMux I__8577 (
            .O(N__35622),
            .I(N__35612));
    InMux I__8576 (
            .O(N__35621),
            .I(N__35608));
    InMux I__8575 (
            .O(N__35620),
            .I(N__35604));
    LocalMux I__8574 (
            .O(N__35617),
            .I(N__35599));
    Span4Mux_h I__8573 (
            .O(N__35612),
            .I(N__35599));
    InMux I__8572 (
            .O(N__35611),
            .I(N__35596));
    LocalMux I__8571 (
            .O(N__35608),
            .I(N__35593));
    InMux I__8570 (
            .O(N__35607),
            .I(N__35590));
    LocalMux I__8569 (
            .O(N__35604),
            .I(N__35585));
    Span4Mux_v I__8568 (
            .O(N__35599),
            .I(N__35585));
    LocalMux I__8567 (
            .O(N__35596),
            .I(N__35582));
    Odrv12 I__8566 (
            .O(N__35593),
            .I(M_this_state_qZ0Z_8));
    LocalMux I__8565 (
            .O(N__35590),
            .I(M_this_state_qZ0Z_8));
    Odrv4 I__8564 (
            .O(N__35585),
            .I(M_this_state_qZ0Z_8));
    Odrv12 I__8563 (
            .O(N__35582),
            .I(M_this_state_qZ0Z_8));
    InMux I__8562 (
            .O(N__35573),
            .I(N__35570));
    LocalMux I__8561 (
            .O(N__35570),
            .I(N__35567));
    Sp12to4 I__8560 (
            .O(N__35567),
            .I(N__35564));
    Span12Mux_v I__8559 (
            .O(N__35564),
            .I(N__35561));
    Odrv12 I__8558 (
            .O(N__35561),
            .I(port_address_in_2));
    InMux I__8557 (
            .O(N__35558),
            .I(N__35555));
    LocalMux I__8556 (
            .O(N__35555),
            .I(N__35552));
    Span4Mux_v I__8555 (
            .O(N__35552),
            .I(N__35549));
    Span4Mux_h I__8554 (
            .O(N__35549),
            .I(N__35546));
    Span4Mux_h I__8553 (
            .O(N__35546),
            .I(N__35543));
    Odrv4 I__8552 (
            .O(N__35543),
            .I(port_address_in_6));
    InMux I__8551 (
            .O(N__35540),
            .I(N__35536));
    InMux I__8550 (
            .O(N__35539),
            .I(N__35533));
    LocalMux I__8549 (
            .O(N__35536),
            .I(N__35530));
    LocalMux I__8548 (
            .O(N__35533),
            .I(N__35527));
    Odrv4 I__8547 (
            .O(N__35530),
            .I(this_vga_signals_M_this_state_d28_0_a2_0_1));
    Odrv4 I__8546 (
            .O(N__35527),
            .I(this_vga_signals_M_this_state_d28_0_a2_0_1));
    CEMux I__8545 (
            .O(N__35522),
            .I(N__35519));
    LocalMux I__8544 (
            .O(N__35519),
            .I(N__35516));
    Span4Mux_h I__8543 (
            .O(N__35516),
            .I(N__35513));
    Span4Mux_h I__8542 (
            .O(N__35513),
            .I(N__35510));
    Odrv4 I__8541 (
            .O(N__35510),
            .I(N_1264_0));
    CascadeMux I__8540 (
            .O(N__35507),
            .I(N__35504));
    InMux I__8539 (
            .O(N__35504),
            .I(N__35500));
    CascadeMux I__8538 (
            .O(N__35503),
            .I(N__35497));
    LocalMux I__8537 (
            .O(N__35500),
            .I(N__35494));
    InMux I__8536 (
            .O(N__35497),
            .I(N__35491));
    Span4Mux_h I__8535 (
            .O(N__35494),
            .I(N__35488));
    LocalMux I__8534 (
            .O(N__35491),
            .I(N__35485));
    Odrv4 I__8533 (
            .O(N__35488),
            .I(\this_start_data_delay.N_387 ));
    Odrv12 I__8532 (
            .O(N__35485),
            .I(\this_start_data_delay.N_387 ));
    InMux I__8531 (
            .O(N__35480),
            .I(N__35477));
    LocalMux I__8530 (
            .O(N__35477),
            .I(N__35473));
    InMux I__8529 (
            .O(N__35476),
            .I(N__35470));
    Span4Mux_h I__8528 (
            .O(N__35473),
            .I(N__35464));
    LocalMux I__8527 (
            .O(N__35470),
            .I(N__35464));
    InMux I__8526 (
            .O(N__35469),
            .I(N__35461));
    Span4Mux_v I__8525 (
            .O(N__35464),
            .I(N__35454));
    LocalMux I__8524 (
            .O(N__35461),
            .I(N__35454));
    InMux I__8523 (
            .O(N__35460),
            .I(N__35451));
    InMux I__8522 (
            .O(N__35459),
            .I(N__35448));
    Span4Mux_v I__8521 (
            .O(N__35454),
            .I(N__35445));
    LocalMux I__8520 (
            .O(N__35451),
            .I(N__35440));
    LocalMux I__8519 (
            .O(N__35448),
            .I(N__35440));
    Span4Mux_v I__8518 (
            .O(N__35445),
            .I(N__35437));
    Span12Mux_h I__8517 (
            .O(N__35440),
            .I(N__35434));
    IoSpan4Mux I__8516 (
            .O(N__35437),
            .I(N__35431));
    Odrv12 I__8515 (
            .O(N__35434),
            .I(port_address_in_0));
    Odrv4 I__8514 (
            .O(N__35431),
            .I(port_address_in_0));
    InMux I__8513 (
            .O(N__35426),
            .I(N__35421));
    InMux I__8512 (
            .O(N__35425),
            .I(N__35418));
    CascadeMux I__8511 (
            .O(N__35424),
            .I(N__35414));
    LocalMux I__8510 (
            .O(N__35421),
            .I(N__35410));
    LocalMux I__8509 (
            .O(N__35418),
            .I(N__35407));
    InMux I__8508 (
            .O(N__35417),
            .I(N__35404));
    InMux I__8507 (
            .O(N__35414),
            .I(N__35401));
    InMux I__8506 (
            .O(N__35413),
            .I(N__35398));
    Span4Mux_v I__8505 (
            .O(N__35410),
            .I(N__35395));
    Span4Mux_h I__8504 (
            .O(N__35407),
            .I(N__35386));
    LocalMux I__8503 (
            .O(N__35404),
            .I(N__35386));
    LocalMux I__8502 (
            .O(N__35401),
            .I(N__35386));
    LocalMux I__8501 (
            .O(N__35398),
            .I(N__35386));
    Sp12to4 I__8500 (
            .O(N__35395),
            .I(N__35383));
    Span4Mux_v I__8499 (
            .O(N__35386),
            .I(N__35380));
    Span12Mux_h I__8498 (
            .O(N__35383),
            .I(N__35377));
    Sp12to4 I__8497 (
            .O(N__35380),
            .I(N__35374));
    Odrv12 I__8496 (
            .O(N__35377),
            .I(port_address_in_4));
    Odrv12 I__8495 (
            .O(N__35374),
            .I(port_address_in_4));
    CascadeMux I__8494 (
            .O(N__35369),
            .I(\this_start_data_delay.N_337_cascade_ ));
    InMux I__8493 (
            .O(N__35366),
            .I(N__35360));
    InMux I__8492 (
            .O(N__35365),
            .I(N__35355));
    InMux I__8491 (
            .O(N__35364),
            .I(N__35355));
    InMux I__8490 (
            .O(N__35363),
            .I(N__35352));
    LocalMux I__8489 (
            .O(N__35360),
            .I(\this_start_data_delay.N_386 ));
    LocalMux I__8488 (
            .O(N__35355),
            .I(\this_start_data_delay.N_386 ));
    LocalMux I__8487 (
            .O(N__35352),
            .I(\this_start_data_delay.N_386 ));
    InMux I__8486 (
            .O(N__35345),
            .I(N__35337));
    InMux I__8485 (
            .O(N__35344),
            .I(N__35337));
    InMux I__8484 (
            .O(N__35343),
            .I(N__35331));
    InMux I__8483 (
            .O(N__35342),
            .I(N__35331));
    LocalMux I__8482 (
            .O(N__35337),
            .I(N__35328));
    InMux I__8481 (
            .O(N__35336),
            .I(N__35325));
    LocalMux I__8480 (
            .O(N__35331),
            .I(N__35322));
    Odrv12 I__8479 (
            .O(N__35328),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    LocalMux I__8478 (
            .O(N__35325),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    Odrv4 I__8477 (
            .O(N__35322),
            .I(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ));
    CascadeMux I__8476 (
            .O(N__35315),
            .I(N__35308));
    InMux I__8475 (
            .O(N__35314),
            .I(N__35303));
    InMux I__8474 (
            .O(N__35313),
            .I(N__35298));
    InMux I__8473 (
            .O(N__35312),
            .I(N__35298));
    InMux I__8472 (
            .O(N__35311),
            .I(N__35295));
    InMux I__8471 (
            .O(N__35308),
            .I(N__35292));
    InMux I__8470 (
            .O(N__35307),
            .I(N__35287));
    InMux I__8469 (
            .O(N__35306),
            .I(N__35287));
    LocalMux I__8468 (
            .O(N__35303),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__8467 (
            .O(N__35298),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__8466 (
            .O(N__35295),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__8465 (
            .O(N__35292),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    LocalMux I__8464 (
            .O(N__35287),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ));
    InMux I__8463 (
            .O(N__35276),
            .I(N__35273));
    LocalMux I__8462 (
            .O(N__35273),
            .I(N__35268));
    InMux I__8461 (
            .O(N__35272),
            .I(N__35264));
    InMux I__8460 (
            .O(N__35271),
            .I(N__35261));
    Span4Mux_h I__8459 (
            .O(N__35268),
            .I(N__35258));
    InMux I__8458 (
            .O(N__35267),
            .I(N__35254));
    LocalMux I__8457 (
            .O(N__35264),
            .I(N__35246));
    LocalMux I__8456 (
            .O(N__35261),
            .I(N__35246));
    Span4Mux_h I__8455 (
            .O(N__35258),
            .I(N__35243));
    InMux I__8454 (
            .O(N__35257),
            .I(N__35240));
    LocalMux I__8453 (
            .O(N__35254),
            .I(N__35236));
    InMux I__8452 (
            .O(N__35253),
            .I(N__35231));
    InMux I__8451 (
            .O(N__35252),
            .I(N__35231));
    CascadeMux I__8450 (
            .O(N__35251),
            .I(N__35227));
    Span12Mux_h I__8449 (
            .O(N__35246),
            .I(N__35224));
    Span4Mux_h I__8448 (
            .O(N__35243),
            .I(N__35221));
    LocalMux I__8447 (
            .O(N__35240),
            .I(N__35218));
    InMux I__8446 (
            .O(N__35239),
            .I(N__35215));
    Span4Mux_v I__8445 (
            .O(N__35236),
            .I(N__35210));
    LocalMux I__8444 (
            .O(N__35231),
            .I(N__35210));
    InMux I__8443 (
            .O(N__35230),
            .I(N__35207));
    InMux I__8442 (
            .O(N__35227),
            .I(N__35204));
    Odrv12 I__8441 (
            .O(N__35224),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__8440 (
            .O(N__35221),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv12 I__8439 (
            .O(N__35218),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__8438 (
            .O(N__35215),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    Odrv4 I__8437 (
            .O(N__35210),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__8436 (
            .O(N__35207),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    LocalMux I__8435 (
            .O(N__35204),
            .I(\this_vga_signals.M_vcounter_qZ0Z_9 ));
    CascadeMux I__8434 (
            .O(N__35189),
            .I(N__35186));
    InMux I__8433 (
            .O(N__35186),
            .I(N__35177));
    InMux I__8432 (
            .O(N__35185),
            .I(N__35174));
    InMux I__8431 (
            .O(N__35184),
            .I(N__35169));
    InMux I__8430 (
            .O(N__35183),
            .I(N__35169));
    InMux I__8429 (
            .O(N__35182),
            .I(N__35164));
    InMux I__8428 (
            .O(N__35181),
            .I(N__35164));
    InMux I__8427 (
            .O(N__35180),
            .I(N__35161));
    LocalMux I__8426 (
            .O(N__35177),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__8425 (
            .O(N__35174),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__8424 (
            .O(N__35169),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__8423 (
            .O(N__35164),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    LocalMux I__8422 (
            .O(N__35161),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ));
    InMux I__8421 (
            .O(N__35150),
            .I(N__35147));
    LocalMux I__8420 (
            .O(N__35147),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_1 ));
    InMux I__8419 (
            .O(N__35144),
            .I(N__35141));
    LocalMux I__8418 (
            .O(N__35141),
            .I(N__35138));
    Odrv4 I__8417 (
            .O(N__35138),
            .I(\this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3 ));
    InMux I__8416 (
            .O(N__35135),
            .I(N__35132));
    LocalMux I__8415 (
            .O(N__35132),
            .I(N__35127));
    InMux I__8414 (
            .O(N__35131),
            .I(N__35124));
    InMux I__8413 (
            .O(N__35130),
            .I(N__35121));
    Span4Mux_v I__8412 (
            .O(N__35127),
            .I(N__35117));
    LocalMux I__8411 (
            .O(N__35124),
            .I(N__35112));
    LocalMux I__8410 (
            .O(N__35121),
            .I(N__35112));
    InMux I__8409 (
            .O(N__35120),
            .I(N__35109));
    Odrv4 I__8408 (
            .O(N__35117),
            .I(\this_start_data_delay.N_424 ));
    Odrv12 I__8407 (
            .O(N__35112),
            .I(\this_start_data_delay.N_424 ));
    LocalMux I__8406 (
            .O(N__35109),
            .I(\this_start_data_delay.N_424 ));
    InMux I__8405 (
            .O(N__35102),
            .I(N__35099));
    LocalMux I__8404 (
            .O(N__35099),
            .I(N__35093));
    InMux I__8403 (
            .O(N__35098),
            .I(N__35090));
    InMux I__8402 (
            .O(N__35097),
            .I(N__35086));
    InMux I__8401 (
            .O(N__35096),
            .I(N__35082));
    Span4Mux_h I__8400 (
            .O(N__35093),
            .I(N__35079));
    LocalMux I__8399 (
            .O(N__35090),
            .I(N__35076));
    InMux I__8398 (
            .O(N__35089),
            .I(N__35073));
    LocalMux I__8397 (
            .O(N__35086),
            .I(N__35069));
    InMux I__8396 (
            .O(N__35085),
            .I(N__35066));
    LocalMux I__8395 (
            .O(N__35082),
            .I(N__35063));
    Span4Mux_v I__8394 (
            .O(N__35079),
            .I(N__35058));
    Span4Mux_h I__8393 (
            .O(N__35076),
            .I(N__35058));
    LocalMux I__8392 (
            .O(N__35073),
            .I(N__35055));
    InMux I__8391 (
            .O(N__35072),
            .I(N__35052));
    Span12Mux_s6_v I__8390 (
            .O(N__35069),
            .I(N__35048));
    LocalMux I__8389 (
            .O(N__35066),
            .I(N__35045));
    Span4Mux_h I__8388 (
            .O(N__35063),
            .I(N__35042));
    Span4Mux_v I__8387 (
            .O(N__35058),
            .I(N__35037));
    Span4Mux_h I__8386 (
            .O(N__35055),
            .I(N__35037));
    LocalMux I__8385 (
            .O(N__35052),
            .I(N__35034));
    InMux I__8384 (
            .O(N__35051),
            .I(N__35031));
    Span12Mux_h I__8383 (
            .O(N__35048),
            .I(N__35028));
    Span12Mux_v I__8382 (
            .O(N__35045),
            .I(N__35025));
    Sp12to4 I__8381 (
            .O(N__35042),
            .I(N__35022));
    Span4Mux_v I__8380 (
            .O(N__35037),
            .I(N__35017));
    Span4Mux_h I__8379 (
            .O(N__35034),
            .I(N__35017));
    LocalMux I__8378 (
            .O(N__35031),
            .I(N__35014));
    Span12Mux_v I__8377 (
            .O(N__35028),
            .I(N__35009));
    Span12Mux_h I__8376 (
            .O(N__35025),
            .I(N__35009));
    Span12Mux_v I__8375 (
            .O(N__35022),
            .I(N__35006));
    Span4Mux_v I__8374 (
            .O(N__35017),
            .I(N__35001));
    Span4Mux_h I__8373 (
            .O(N__35014),
            .I(N__35001));
    Odrv12 I__8372 (
            .O(N__35009),
            .I(M_this_spr_ram_write_data_0));
    Odrv12 I__8371 (
            .O(N__35006),
            .I(M_this_spr_ram_write_data_0));
    Odrv4 I__8370 (
            .O(N__35001),
            .I(M_this_spr_ram_write_data_0));
    InMux I__8369 (
            .O(N__34994),
            .I(N__34990));
    InMux I__8368 (
            .O(N__34993),
            .I(N__34987));
    LocalMux I__8367 (
            .O(N__34990),
            .I(N__34981));
    LocalMux I__8366 (
            .O(N__34987),
            .I(N__34978));
    InMux I__8365 (
            .O(N__34986),
            .I(N__34975));
    InMux I__8364 (
            .O(N__34985),
            .I(N__34970));
    InMux I__8363 (
            .O(N__34984),
            .I(N__34967));
    Span12Mux_h I__8362 (
            .O(N__34981),
            .I(N__34964));
    Span4Mux_h I__8361 (
            .O(N__34978),
            .I(N__34959));
    LocalMux I__8360 (
            .O(N__34975),
            .I(N__34959));
    InMux I__8359 (
            .O(N__34974),
            .I(N__34954));
    InMux I__8358 (
            .O(N__34973),
            .I(N__34954));
    LocalMux I__8357 (
            .O(N__34970),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__8356 (
            .O(N__34967),
            .I(M_this_state_qZ0Z_11));
    Odrv12 I__8355 (
            .O(N__34964),
            .I(M_this_state_qZ0Z_11));
    Odrv4 I__8354 (
            .O(N__34959),
            .I(M_this_state_qZ0Z_11));
    LocalMux I__8353 (
            .O(N__34954),
            .I(M_this_state_qZ0Z_11));
    CascadeMux I__8352 (
            .O(N__34943),
            .I(\this_start_data_delay.N_245_0_cascade_ ));
    InMux I__8351 (
            .O(N__34940),
            .I(N__34937));
    LocalMux I__8350 (
            .O(N__34937),
            .I(N__34934));
    Odrv12 I__8349 (
            .O(N__34934),
            .I(un20_i_a4_0_a2_0_a2_1));
    InMux I__8348 (
            .O(N__34931),
            .I(N__34927));
    InMux I__8347 (
            .O(N__34930),
            .I(N__34923));
    LocalMux I__8346 (
            .O(N__34927),
            .I(N__34920));
    InMux I__8345 (
            .O(N__34926),
            .I(N__34917));
    LocalMux I__8344 (
            .O(N__34923),
            .I(N__34913));
    Span4Mux_v I__8343 (
            .O(N__34920),
            .I(N__34908));
    LocalMux I__8342 (
            .O(N__34917),
            .I(N__34908));
    CascadeMux I__8341 (
            .O(N__34916),
            .I(N__34904));
    Span4Mux_v I__8340 (
            .O(N__34913),
            .I(N__34898));
    Span4Mux_h I__8339 (
            .O(N__34908),
            .I(N__34898));
    CascadeMux I__8338 (
            .O(N__34907),
            .I(N__34895));
    InMux I__8337 (
            .O(N__34904),
            .I(N__34889));
    InMux I__8336 (
            .O(N__34903),
            .I(N__34886));
    Span4Mux_h I__8335 (
            .O(N__34898),
            .I(N__34883));
    InMux I__8334 (
            .O(N__34895),
            .I(N__34880));
    CascadeMux I__8333 (
            .O(N__34894),
            .I(N__34877));
    InMux I__8332 (
            .O(N__34893),
            .I(N__34872));
    InMux I__8331 (
            .O(N__34892),
            .I(N__34872));
    LocalMux I__8330 (
            .O(N__34889),
            .I(N__34869));
    LocalMux I__8329 (
            .O(N__34886),
            .I(N__34862));
    Span4Mux_v I__8328 (
            .O(N__34883),
            .I(N__34862));
    LocalMux I__8327 (
            .O(N__34880),
            .I(N__34862));
    InMux I__8326 (
            .O(N__34877),
            .I(N__34859));
    LocalMux I__8325 (
            .O(N__34872),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8324 (
            .O(N__34869),
            .I(M_this_state_qZ0Z_13));
    Odrv4 I__8323 (
            .O(N__34862),
            .I(M_this_state_qZ0Z_13));
    LocalMux I__8322 (
            .O(N__34859),
            .I(M_this_state_qZ0Z_13));
    InMux I__8321 (
            .O(N__34850),
            .I(N__34847));
    LocalMux I__8320 (
            .O(N__34847),
            .I(N__34844));
    Odrv12 I__8319 (
            .O(N__34844),
            .I(un20_i_a4_0_a2_2));
    InMux I__8318 (
            .O(N__34841),
            .I(N__34838));
    LocalMux I__8317 (
            .O(N__34838),
            .I(N__34824));
    InMux I__8316 (
            .O(N__34837),
            .I(N__34819));
    InMux I__8315 (
            .O(N__34836),
            .I(N__34819));
    InMux I__8314 (
            .O(N__34835),
            .I(N__34814));
    InMux I__8313 (
            .O(N__34834),
            .I(N__34814));
    InMux I__8312 (
            .O(N__34833),
            .I(N__34805));
    InMux I__8311 (
            .O(N__34832),
            .I(N__34805));
    InMux I__8310 (
            .O(N__34831),
            .I(N__34805));
    InMux I__8309 (
            .O(N__34830),
            .I(N__34805));
    InMux I__8308 (
            .O(N__34829),
            .I(N__34800));
    InMux I__8307 (
            .O(N__34828),
            .I(N__34800));
    InMux I__8306 (
            .O(N__34827),
            .I(N__34797));
    Odrv4 I__8305 (
            .O(N__34824),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__8304 (
            .O(N__34819),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__8303 (
            .O(N__34814),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__8302 (
            .O(N__34805),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__8301 (
            .O(N__34800),
            .I(\this_vga_signals.vaddress_c2 ));
    LocalMux I__8300 (
            .O(N__34797),
            .I(\this_vga_signals.vaddress_c2 ));
    CascadeMux I__8299 (
            .O(N__34784),
            .I(N__34781));
    InMux I__8298 (
            .O(N__34781),
            .I(N__34778));
    LocalMux I__8297 (
            .O(N__34778),
            .I(\this_vga_signals.N_13 ));
    InMux I__8296 (
            .O(N__34775),
            .I(N__34772));
    LocalMux I__8295 (
            .O(N__34772),
            .I(N__34768));
    InMux I__8294 (
            .O(N__34771),
            .I(N__34765));
    Span4Mux_h I__8293 (
            .O(N__34768),
            .I(N__34760));
    LocalMux I__8292 (
            .O(N__34765),
            .I(N__34760));
    Span4Mux_h I__8291 (
            .O(N__34760),
            .I(N__34757));
    Odrv4 I__8290 (
            .O(N__34757),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ));
    InMux I__8289 (
            .O(N__34754),
            .I(N__34749));
    CascadeMux I__8288 (
            .O(N__34753),
            .I(N__34746));
    InMux I__8287 (
            .O(N__34752),
            .I(N__34742));
    LocalMux I__8286 (
            .O(N__34749),
            .I(N__34739));
    InMux I__8285 (
            .O(N__34746),
            .I(N__34734));
    InMux I__8284 (
            .O(N__34745),
            .I(N__34734));
    LocalMux I__8283 (
            .O(N__34742),
            .I(N__34725));
    Span4Mux_h I__8282 (
            .O(N__34739),
            .I(N__34720));
    LocalMux I__8281 (
            .O(N__34734),
            .I(N__34720));
    InMux I__8280 (
            .O(N__34733),
            .I(N__34717));
    InMux I__8279 (
            .O(N__34732),
            .I(N__34713));
    InMux I__8278 (
            .O(N__34731),
            .I(N__34708));
    InMux I__8277 (
            .O(N__34730),
            .I(N__34708));
    InMux I__8276 (
            .O(N__34729),
            .I(N__34703));
    InMux I__8275 (
            .O(N__34728),
            .I(N__34703));
    Span4Mux_h I__8274 (
            .O(N__34725),
            .I(N__34696));
    Span4Mux_v I__8273 (
            .O(N__34720),
            .I(N__34696));
    LocalMux I__8272 (
            .O(N__34717),
            .I(N__34696));
    InMux I__8271 (
            .O(N__34716),
            .I(N__34693));
    LocalMux I__8270 (
            .O(N__34713),
            .I(N__34686));
    LocalMux I__8269 (
            .O(N__34708),
            .I(N__34686));
    LocalMux I__8268 (
            .O(N__34703),
            .I(N__34686));
    Span4Mux_h I__8267 (
            .O(N__34696),
            .I(N__34683));
    LocalMux I__8266 (
            .O(N__34693),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv12 I__8265 (
            .O(N__34686),
            .I(this_vga_signals_M_vcounter_q_7));
    Odrv4 I__8264 (
            .O(N__34683),
            .I(this_vga_signals_M_vcounter_q_7));
    InMux I__8263 (
            .O(N__34676),
            .I(N__34673));
    LocalMux I__8262 (
            .O(N__34673),
            .I(N__34669));
    InMux I__8261 (
            .O(N__34672),
            .I(N__34666));
    Span4Mux_h I__8260 (
            .O(N__34669),
            .I(N__34661));
    LocalMux I__8259 (
            .O(N__34666),
            .I(N__34661));
    Span4Mux_h I__8258 (
            .O(N__34661),
            .I(N__34658));
    Odrv4 I__8257 (
            .O(N__34658),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ));
    CascadeMux I__8256 (
            .O(N__34655),
            .I(N__34652));
    InMux I__8255 (
            .O(N__34652),
            .I(N__34644));
    InMux I__8254 (
            .O(N__34651),
            .I(N__34644));
    InMux I__8253 (
            .O(N__34650),
            .I(N__34641));
    InMux I__8252 (
            .O(N__34649),
            .I(N__34637));
    LocalMux I__8251 (
            .O(N__34644),
            .I(N__34634));
    LocalMux I__8250 (
            .O(N__34641),
            .I(N__34629));
    CascadeMux I__8249 (
            .O(N__34640),
            .I(N__34623));
    LocalMux I__8248 (
            .O(N__34637),
            .I(N__34617));
    Span4Mux_h I__8247 (
            .O(N__34634),
            .I(N__34617));
    InMux I__8246 (
            .O(N__34633),
            .I(N__34614));
    CascadeMux I__8245 (
            .O(N__34632),
            .I(N__34611));
    Span4Mux_v I__8244 (
            .O(N__34629),
            .I(N__34608));
    InMux I__8243 (
            .O(N__34628),
            .I(N__34605));
    InMux I__8242 (
            .O(N__34627),
            .I(N__34600));
    InMux I__8241 (
            .O(N__34626),
            .I(N__34600));
    InMux I__8240 (
            .O(N__34623),
            .I(N__34595));
    InMux I__8239 (
            .O(N__34622),
            .I(N__34595));
    Span4Mux_h I__8238 (
            .O(N__34617),
            .I(N__34592));
    LocalMux I__8237 (
            .O(N__34614),
            .I(N__34589));
    InMux I__8236 (
            .O(N__34611),
            .I(N__34586));
    Span4Mux_h I__8235 (
            .O(N__34608),
            .I(N__34577));
    LocalMux I__8234 (
            .O(N__34605),
            .I(N__34577));
    LocalMux I__8233 (
            .O(N__34600),
            .I(N__34577));
    LocalMux I__8232 (
            .O(N__34595),
            .I(N__34577));
    Odrv4 I__8231 (
            .O(N__34592),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv12 I__8230 (
            .O(N__34589),
            .I(this_vga_signals_M_vcounter_q_8));
    LocalMux I__8229 (
            .O(N__34586),
            .I(this_vga_signals_M_vcounter_q_8));
    Odrv4 I__8228 (
            .O(N__34577),
            .I(this_vga_signals_M_vcounter_q_8));
    InMux I__8227 (
            .O(N__34568),
            .I(N__34565));
    LocalMux I__8226 (
            .O(N__34565),
            .I(N__34561));
    InMux I__8225 (
            .O(N__34564),
            .I(N__34558));
    Span4Mux_v I__8224 (
            .O(N__34561),
            .I(N__34553));
    LocalMux I__8223 (
            .O(N__34558),
            .I(N__34553));
    Span4Mux_h I__8222 (
            .O(N__34553),
            .I(N__34550));
    Odrv4 I__8221 (
            .O(N__34550),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ));
    InMux I__8220 (
            .O(N__34547),
            .I(N__34543));
    InMux I__8219 (
            .O(N__34546),
            .I(N__34540));
    LocalMux I__8218 (
            .O(N__34543),
            .I(N__34536));
    LocalMux I__8217 (
            .O(N__34540),
            .I(N__34533));
    InMux I__8216 (
            .O(N__34539),
            .I(N__34530));
    Span4Mux_h I__8215 (
            .O(N__34536),
            .I(N__34527));
    Span4Mux_v I__8214 (
            .O(N__34533),
            .I(N__34522));
    LocalMux I__8213 (
            .O(N__34530),
            .I(N__34522));
    Span4Mux_h I__8212 (
            .O(N__34527),
            .I(N__34519));
    Span4Mux_h I__8211 (
            .O(N__34522),
            .I(N__34516));
    Odrv4 I__8210 (
            .O(N__34519),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    Odrv4 I__8209 (
            .O(N__34516),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ));
    CEMux I__8208 (
            .O(N__34511),
            .I(N__34505));
    CEMux I__8207 (
            .O(N__34510),
            .I(N__34502));
    CEMux I__8206 (
            .O(N__34509),
            .I(N__34499));
    CEMux I__8205 (
            .O(N__34508),
            .I(N__34495));
    LocalMux I__8204 (
            .O(N__34505),
            .I(N__34492));
    LocalMux I__8203 (
            .O(N__34502),
            .I(N__34488));
    LocalMux I__8202 (
            .O(N__34499),
            .I(N__34485));
    CEMux I__8201 (
            .O(N__34498),
            .I(N__34481));
    LocalMux I__8200 (
            .O(N__34495),
            .I(N__34476));
    Span4Mux_v I__8199 (
            .O(N__34492),
            .I(N__34476));
    CEMux I__8198 (
            .O(N__34491),
            .I(N__34473));
    Span4Mux_v I__8197 (
            .O(N__34488),
            .I(N__34468));
    Span4Mux_v I__8196 (
            .O(N__34485),
            .I(N__34468));
    CEMux I__8195 (
            .O(N__34484),
            .I(N__34465));
    LocalMux I__8194 (
            .O(N__34481),
            .I(N__34462));
    Span4Mux_h I__8193 (
            .O(N__34476),
            .I(N__34459));
    LocalMux I__8192 (
            .O(N__34473),
            .I(N__34454));
    Span4Mux_h I__8191 (
            .O(N__34468),
            .I(N__34454));
    LocalMux I__8190 (
            .O(N__34465),
            .I(N__34451));
    Span4Mux_h I__8189 (
            .O(N__34462),
            .I(N__34448));
    Span4Mux_h I__8188 (
            .O(N__34459),
            .I(N__34445));
    Span4Mux_h I__8187 (
            .O(N__34454),
            .I(N__34442));
    Odrv12 I__8186 (
            .O(N__34451),
            .I(\this_vga_signals.N_933_0 ));
    Odrv4 I__8185 (
            .O(N__34448),
            .I(\this_vga_signals.N_933_0 ));
    Odrv4 I__8184 (
            .O(N__34445),
            .I(\this_vga_signals.N_933_0 ));
    Odrv4 I__8183 (
            .O(N__34442),
            .I(\this_vga_signals.N_933_0 ));
    SRMux I__8182 (
            .O(N__34433),
            .I(N__34409));
    SRMux I__8181 (
            .O(N__34432),
            .I(N__34409));
    SRMux I__8180 (
            .O(N__34431),
            .I(N__34409));
    SRMux I__8179 (
            .O(N__34430),
            .I(N__34409));
    SRMux I__8178 (
            .O(N__34429),
            .I(N__34409));
    SRMux I__8177 (
            .O(N__34428),
            .I(N__34409));
    SRMux I__8176 (
            .O(N__34427),
            .I(N__34409));
    SRMux I__8175 (
            .O(N__34426),
            .I(N__34409));
    GlobalMux I__8174 (
            .O(N__34409),
            .I(N__34406));
    gio2CtrlBuf I__8173 (
            .O(N__34406),
            .I(\this_vga_signals.N_1188_g ));
    CascadeMux I__8172 (
            .O(N__34403),
            .I(N_422_2_cascade_));
    IoInMux I__8171 (
            .O(N__34400),
            .I(N__34397));
    LocalMux I__8170 (
            .O(N__34397),
            .I(N__34394));
    Span4Mux_s0_h I__8169 (
            .O(N__34394),
            .I(N__34391));
    Span4Mux_v I__8168 (
            .O(N__34391),
            .I(N__34388));
    Sp12to4 I__8167 (
            .O(N__34388),
            .I(N__34385));
    Span12Mux_v I__8166 (
            .O(N__34385),
            .I(N__34382));
    Odrv12 I__8165 (
            .O(N__34382),
            .I(N_458_i));
    CascadeMux I__8164 (
            .O(N__34379),
            .I(N__34376));
    InMux I__8163 (
            .O(N__34376),
            .I(N__34373));
    LocalMux I__8162 (
            .O(N__34373),
            .I(\this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6 ));
    InMux I__8161 (
            .O(N__34370),
            .I(N__34362));
    InMux I__8160 (
            .O(N__34369),
            .I(N__34362));
    InMux I__8159 (
            .O(N__34368),
            .I(N__34357));
    InMux I__8158 (
            .O(N__34367),
            .I(N__34357));
    LocalMux I__8157 (
            .O(N__34362),
            .I(M_this_substate_qZ0));
    LocalMux I__8156 (
            .O(N__34357),
            .I(M_this_substate_qZ0));
    InMux I__8155 (
            .O(N__34352),
            .I(N__34345));
    InMux I__8154 (
            .O(N__34351),
            .I(N__34345));
    InMux I__8153 (
            .O(N__34350),
            .I(N__34342));
    LocalMux I__8152 (
            .O(N__34345),
            .I(N__34339));
    LocalMux I__8151 (
            .O(N__34342),
            .I(N__34336));
    Odrv4 I__8150 (
            .O(N__34339),
            .I(\this_start_data_delay.N_467 ));
    Odrv12 I__8149 (
            .O(N__34336),
            .I(\this_start_data_delay.N_467 ));
    CascadeMux I__8148 (
            .O(N__34331),
            .I(\this_start_data_delay.N_386_cascade_ ));
    CascadeMux I__8147 (
            .O(N__34328),
            .I(N__34322));
    InMux I__8146 (
            .O(N__34327),
            .I(N__34319));
    InMux I__8145 (
            .O(N__34326),
            .I(N__34312));
    InMux I__8144 (
            .O(N__34325),
            .I(N__34312));
    InMux I__8143 (
            .O(N__34322),
            .I(N__34312));
    LocalMux I__8142 (
            .O(N__34319),
            .I(N__34307));
    LocalMux I__8141 (
            .O(N__34312),
            .I(N__34307));
    Span12Mux_h I__8140 (
            .O(N__34307),
            .I(N__34304));
    Odrv12 I__8139 (
            .O(N__34304),
            .I(port_address_in_1));
    InMux I__8138 (
            .O(N__34301),
            .I(N__34292));
    InMux I__8137 (
            .O(N__34300),
            .I(N__34292));
    InMux I__8136 (
            .O(N__34299),
            .I(N__34292));
    LocalMux I__8135 (
            .O(N__34292),
            .I(\this_start_data_delay.N_380 ));
    InMux I__8134 (
            .O(N__34289),
            .I(N__34286));
    LocalMux I__8133 (
            .O(N__34286),
            .I(\this_start_data_delay.N_341 ));
    InMux I__8132 (
            .O(N__34283),
            .I(N__34279));
    InMux I__8131 (
            .O(N__34282),
            .I(N__34273));
    LocalMux I__8130 (
            .O(N__34279),
            .I(N__34270));
    InMux I__8129 (
            .O(N__34278),
            .I(N__34267));
    InMux I__8128 (
            .O(N__34277),
            .I(N__34264));
    InMux I__8127 (
            .O(N__34276),
            .I(N__34260));
    LocalMux I__8126 (
            .O(N__34273),
            .I(N__34257));
    Span4Mux_v I__8125 (
            .O(N__34270),
            .I(N__34252));
    LocalMux I__8124 (
            .O(N__34267),
            .I(N__34252));
    LocalMux I__8123 (
            .O(N__34264),
            .I(N__34249));
    InMux I__8122 (
            .O(N__34263),
            .I(N__34246));
    LocalMux I__8121 (
            .O(N__34260),
            .I(N__34241));
    Sp12to4 I__8120 (
            .O(N__34257),
            .I(N__34238));
    Span4Mux_v I__8119 (
            .O(N__34252),
            .I(N__34235));
    Span4Mux_h I__8118 (
            .O(N__34249),
            .I(N__34232));
    LocalMux I__8117 (
            .O(N__34246),
            .I(N__34229));
    InMux I__8116 (
            .O(N__34245),
            .I(N__34226));
    InMux I__8115 (
            .O(N__34244),
            .I(N__34223));
    Span12Mux_s8_h I__8114 (
            .O(N__34241),
            .I(N__34220));
    Span12Mux_v I__8113 (
            .O(N__34238),
            .I(N__34217));
    Sp12to4 I__8112 (
            .O(N__34235),
            .I(N__34214));
    Span4Mux_v I__8111 (
            .O(N__34232),
            .I(N__34209));
    Span4Mux_h I__8110 (
            .O(N__34229),
            .I(N__34209));
    LocalMux I__8109 (
            .O(N__34226),
            .I(N__34206));
    LocalMux I__8108 (
            .O(N__34223),
            .I(N__34203));
    Span12Mux_h I__8107 (
            .O(N__34220),
            .I(N__34200));
    Span12Mux_h I__8106 (
            .O(N__34217),
            .I(N__34195));
    Span12Mux_h I__8105 (
            .O(N__34214),
            .I(N__34195));
    Span4Mux_v I__8104 (
            .O(N__34209),
            .I(N__34188));
    Span4Mux_h I__8103 (
            .O(N__34206),
            .I(N__34188));
    Span4Mux_h I__8102 (
            .O(N__34203),
            .I(N__34188));
    Odrv12 I__8101 (
            .O(N__34200),
            .I(M_this_spr_ram_write_data_2));
    Odrv12 I__8100 (
            .O(N__34195),
            .I(M_this_spr_ram_write_data_2));
    Odrv4 I__8099 (
            .O(N__34188),
            .I(M_this_spr_ram_write_data_2));
    CascadeMux I__8098 (
            .O(N__34181),
            .I(dma_axb0_cascade_));
    InMux I__8097 (
            .O(N__34178),
            .I(N__34174));
    IoInMux I__8096 (
            .O(N__34177),
            .I(N__34170));
    LocalMux I__8095 (
            .O(N__34174),
            .I(N__34167));
    InMux I__8094 (
            .O(N__34173),
            .I(N__34164));
    LocalMux I__8093 (
            .O(N__34170),
            .I(N__34161));
    Span4Mux_v I__8092 (
            .O(N__34167),
            .I(N__34158));
    LocalMux I__8091 (
            .O(N__34164),
            .I(N__34155));
    Span12Mux_s2_h I__8090 (
            .O(N__34161),
            .I(N__34150));
    Sp12to4 I__8089 (
            .O(N__34158),
            .I(N__34147));
    Span4Mux_v I__8088 (
            .O(N__34155),
            .I(N__34144));
    InMux I__8087 (
            .O(N__34154),
            .I(N__34141));
    InMux I__8086 (
            .O(N__34153),
            .I(N__34138));
    Span12Mux_h I__8085 (
            .O(N__34150),
            .I(N__34135));
    Span12Mux_s8_h I__8084 (
            .O(N__34147),
            .I(N__34132));
    Sp12to4 I__8083 (
            .O(N__34144),
            .I(N__34129));
    LocalMux I__8082 (
            .O(N__34141),
            .I(N__34124));
    LocalMux I__8081 (
            .O(N__34138),
            .I(N__34124));
    Span12Mux_v I__8080 (
            .O(N__34135),
            .I(N__34121));
    Span12Mux_h I__8079 (
            .O(N__34132),
            .I(N__34116));
    Span12Mux_h I__8078 (
            .O(N__34129),
            .I(N__34116));
    Span4Mux_h I__8077 (
            .O(N__34124),
            .I(N__34113));
    Odrv12 I__8076 (
            .O(N__34121),
            .I(dma_0));
    Odrv12 I__8075 (
            .O(N__34116),
            .I(dma_0));
    Odrv4 I__8074 (
            .O(N__34113),
            .I(dma_0));
    InMux I__8073 (
            .O(N__34106),
            .I(N__34103));
    LocalMux I__8072 (
            .O(N__34103),
            .I(dma_axb3));
    CascadeMux I__8071 (
            .O(N__34100),
            .I(\this_start_data_delay.N_345_cascade_ ));
    InMux I__8070 (
            .O(N__34097),
            .I(N__34094));
    LocalMux I__8069 (
            .O(N__34094),
            .I(N__34091));
    Odrv12 I__8068 (
            .O(N__34091),
            .I(\this_start_data_delay.N_284_0 ));
    CascadeMux I__8067 (
            .O(N__34088),
            .I(\this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_ ));
    CascadeMux I__8066 (
            .O(N__34085),
            .I(\this_start_data_delay.N_23_1_0_cascade_ ));
    CascadeMux I__8065 (
            .O(N__34082),
            .I(\this_start_data_delay.N_339_cascade_ ));
    CascadeMux I__8064 (
            .O(N__34079),
            .I(\this_vga_signals.m47_0_1_cascade_ ));
    CascadeMux I__8063 (
            .O(N__34076),
            .I(N__34070));
    CascadeMux I__8062 (
            .O(N__34075),
            .I(N__34066));
    CascadeMux I__8061 (
            .O(N__34074),
            .I(N__34062));
    InMux I__8060 (
            .O(N__34073),
            .I(N__34057));
    InMux I__8059 (
            .O(N__34070),
            .I(N__34054));
    InMux I__8058 (
            .O(N__34069),
            .I(N__34049));
    InMux I__8057 (
            .O(N__34066),
            .I(N__34049));
    CascadeMux I__8056 (
            .O(N__34065),
            .I(N__34046));
    InMux I__8055 (
            .O(N__34062),
            .I(N__34042));
    InMux I__8054 (
            .O(N__34061),
            .I(N__34038));
    InMux I__8053 (
            .O(N__34060),
            .I(N__34035));
    LocalMux I__8052 (
            .O(N__34057),
            .I(N__34032));
    LocalMux I__8051 (
            .O(N__34054),
            .I(N__34029));
    LocalMux I__8050 (
            .O(N__34049),
            .I(N__34026));
    InMux I__8049 (
            .O(N__34046),
            .I(N__34023));
    InMux I__8048 (
            .O(N__34045),
            .I(N__34020));
    LocalMux I__8047 (
            .O(N__34042),
            .I(N__34013));
    InMux I__8046 (
            .O(N__34041),
            .I(N__34009));
    LocalMux I__8045 (
            .O(N__34038),
            .I(N__34006));
    LocalMux I__8044 (
            .O(N__34035),
            .I(N__34001));
    Span4Mux_v I__8043 (
            .O(N__34032),
            .I(N__34001));
    Span4Mux_h I__8042 (
            .O(N__34029),
            .I(N__33992));
    Span4Mux_v I__8041 (
            .O(N__34026),
            .I(N__33992));
    LocalMux I__8040 (
            .O(N__34023),
            .I(N__33992));
    LocalMux I__8039 (
            .O(N__34020),
            .I(N__33992));
    InMux I__8038 (
            .O(N__34019),
            .I(N__33987));
    InMux I__8037 (
            .O(N__34018),
            .I(N__33987));
    CascadeMux I__8036 (
            .O(N__34017),
            .I(N__33984));
    CascadeMux I__8035 (
            .O(N__34016),
            .I(N__33981));
    Span4Mux_v I__8034 (
            .O(N__34013),
            .I(N__33977));
    InMux I__8033 (
            .O(N__34012),
            .I(N__33974));
    LocalMux I__8032 (
            .O(N__34009),
            .I(N__33965));
    Span4Mux_v I__8031 (
            .O(N__34006),
            .I(N__33965));
    Span4Mux_h I__8030 (
            .O(N__34001),
            .I(N__33965));
    Span4Mux_v I__8029 (
            .O(N__33992),
            .I(N__33965));
    LocalMux I__8028 (
            .O(N__33987),
            .I(N__33962));
    InMux I__8027 (
            .O(N__33984),
            .I(N__33955));
    InMux I__8026 (
            .O(N__33981),
            .I(N__33955));
    InMux I__8025 (
            .O(N__33980),
            .I(N__33955));
    Odrv4 I__8024 (
            .O(N__33977),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__8023 (
            .O(N__33974),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__8022 (
            .O(N__33965),
            .I(this_vga_signals_M_vcounter_q_6));
    Odrv4 I__8021 (
            .O(N__33962),
            .I(this_vga_signals_M_vcounter_q_6));
    LocalMux I__8020 (
            .O(N__33955),
            .I(this_vga_signals_M_vcounter_q_6));
    CascadeMux I__8019 (
            .O(N__33944),
            .I(N__33935));
    CascadeMux I__8018 (
            .O(N__33943),
            .I(N__33932));
    InMux I__8017 (
            .O(N__33942),
            .I(N__33922));
    InMux I__8016 (
            .O(N__33941),
            .I(N__33919));
    InMux I__8015 (
            .O(N__33940),
            .I(N__33916));
    InMux I__8014 (
            .O(N__33939),
            .I(N__33913));
    InMux I__8013 (
            .O(N__33938),
            .I(N__33908));
    InMux I__8012 (
            .O(N__33935),
            .I(N__33908));
    InMux I__8011 (
            .O(N__33932),
            .I(N__33904));
    InMux I__8010 (
            .O(N__33931),
            .I(N__33898));
    InMux I__8009 (
            .O(N__33930),
            .I(N__33895));
    InMux I__8008 (
            .O(N__33929),
            .I(N__33890));
    InMux I__8007 (
            .O(N__33928),
            .I(N__33890));
    CascadeMux I__8006 (
            .O(N__33927),
            .I(N__33887));
    InMux I__8005 (
            .O(N__33926),
            .I(N__33884));
    InMux I__8004 (
            .O(N__33925),
            .I(N__33881));
    LocalMux I__8003 (
            .O(N__33922),
            .I(N__33878));
    LocalMux I__8002 (
            .O(N__33919),
            .I(N__33868));
    LocalMux I__8001 (
            .O(N__33916),
            .I(N__33868));
    LocalMux I__8000 (
            .O(N__33913),
            .I(N__33865));
    LocalMux I__7999 (
            .O(N__33908),
            .I(N__33862));
    InMux I__7998 (
            .O(N__33907),
            .I(N__33859));
    LocalMux I__7997 (
            .O(N__33904),
            .I(N__33856));
    InMux I__7996 (
            .O(N__33903),
            .I(N__33851));
    InMux I__7995 (
            .O(N__33902),
            .I(N__33851));
    InMux I__7994 (
            .O(N__33901),
            .I(N__33848));
    LocalMux I__7993 (
            .O(N__33898),
            .I(N__33841));
    LocalMux I__7992 (
            .O(N__33895),
            .I(N__33841));
    LocalMux I__7991 (
            .O(N__33890),
            .I(N__33841));
    InMux I__7990 (
            .O(N__33887),
            .I(N__33838));
    LocalMux I__7989 (
            .O(N__33884),
            .I(N__33835));
    LocalMux I__7988 (
            .O(N__33881),
            .I(N__33830));
    Span4Mux_h I__7987 (
            .O(N__33878),
            .I(N__33830));
    InMux I__7986 (
            .O(N__33877),
            .I(N__33823));
    InMux I__7985 (
            .O(N__33876),
            .I(N__33823));
    InMux I__7984 (
            .O(N__33875),
            .I(N__33823));
    InMux I__7983 (
            .O(N__33874),
            .I(N__33818));
    InMux I__7982 (
            .O(N__33873),
            .I(N__33818));
    Span4Mux_v I__7981 (
            .O(N__33868),
            .I(N__33807));
    Span4Mux_v I__7980 (
            .O(N__33865),
            .I(N__33807));
    Span4Mux_v I__7979 (
            .O(N__33862),
            .I(N__33807));
    LocalMux I__7978 (
            .O(N__33859),
            .I(N__33807));
    Span4Mux_v I__7977 (
            .O(N__33856),
            .I(N__33807));
    LocalMux I__7976 (
            .O(N__33851),
            .I(N__33802));
    LocalMux I__7975 (
            .O(N__33848),
            .I(N__33802));
    Odrv4 I__7974 (
            .O(N__33841),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__7973 (
            .O(N__33838),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__7972 (
            .O(N__33835),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__7971 (
            .O(N__33830),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__7970 (
            .O(N__33823),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    LocalMux I__7969 (
            .O(N__33818),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv4 I__7968 (
            .O(N__33807),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    Odrv12 I__7967 (
            .O(N__33802),
            .I(\this_vga_signals.M_vcounter_qZ0Z_4 ));
    CascadeMux I__7966 (
            .O(N__33785),
            .I(\this_vga_signals.SUM_2_cascade_ ));
    InMux I__7965 (
            .O(N__33782),
            .I(N__33779));
    LocalMux I__7964 (
            .O(N__33779),
            .I(\this_vga_signals.g0_0_i_a7_1 ));
    CascadeMux I__7963 (
            .O(N__33776),
            .I(N__33773));
    InMux I__7962 (
            .O(N__33773),
            .I(N__33770));
    LocalMux I__7961 (
            .O(N__33770),
            .I(N__33767));
    Odrv4 I__7960 (
            .O(N__33767),
            .I(N_88));
    InMux I__7959 (
            .O(N__33764),
            .I(N__33758));
    InMux I__7958 (
            .O(N__33763),
            .I(N__33758));
    LocalMux I__7957 (
            .O(N__33758),
            .I(N__33755));
    Span12Mux_v I__7956 (
            .O(N__33755),
            .I(N__33752));
    Span12Mux_h I__7955 (
            .O(N__33752),
            .I(N__33749));
    Odrv12 I__7954 (
            .O(N__33749),
            .I(port_address_in_5));
    CascadeMux I__7953 (
            .O(N__33746),
            .I(N__33743));
    InMux I__7952 (
            .O(N__33743),
            .I(N__33737));
    InMux I__7951 (
            .O(N__33742),
            .I(N__33737));
    LocalMux I__7950 (
            .O(N__33737),
            .I(N__33734));
    Span4Mux_v I__7949 (
            .O(N__33734),
            .I(N__33731));
    Sp12to4 I__7948 (
            .O(N__33731),
            .I(N__33728));
    Span12Mux_h I__7947 (
            .O(N__33728),
            .I(N__33725));
    Span12Mux_v I__7946 (
            .O(N__33725),
            .I(N__33722));
    Odrv12 I__7945 (
            .O(N__33722),
            .I(port_address_in_7));
    InMux I__7944 (
            .O(N__33719),
            .I(N__33713));
    InMux I__7943 (
            .O(N__33718),
            .I(N__33713));
    LocalMux I__7942 (
            .O(N__33713),
            .I(N__33710));
    Span12Mux_v I__7941 (
            .O(N__33710),
            .I(N__33707));
    Span12Mux_h I__7940 (
            .O(N__33707),
            .I(N__33704));
    Odrv12 I__7939 (
            .O(N__33704),
            .I(port_address_in_3));
    CascadeMux I__7938 (
            .O(N__33701),
            .I(N__33698));
    InMux I__7937 (
            .O(N__33698),
            .I(N__33695));
    LocalMux I__7936 (
            .O(N__33695),
            .I(N__33692));
    Odrv4 I__7935 (
            .O(N__33692),
            .I(\this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6 ));
    InMux I__7934 (
            .O(N__33689),
            .I(N__33684));
    InMux I__7933 (
            .O(N__33688),
            .I(N__33681));
    InMux I__7932 (
            .O(N__33687),
            .I(N__33678));
    LocalMux I__7931 (
            .O(N__33684),
            .I(N__33673));
    LocalMux I__7930 (
            .O(N__33681),
            .I(N__33673));
    LocalMux I__7929 (
            .O(N__33678),
            .I(N__33670));
    Span4Mux_v I__7928 (
            .O(N__33673),
            .I(N__33667));
    Span4Mux_h I__7927 (
            .O(N__33670),
            .I(N__33664));
    Odrv4 I__7926 (
            .O(N__33667),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    Odrv4 I__7925 (
            .O(N__33664),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ));
    InMux I__7924 (
            .O(N__33659),
            .I(N__33653));
    InMux I__7923 (
            .O(N__33658),
            .I(N__33646));
    InMux I__7922 (
            .O(N__33657),
            .I(N__33646));
    InMux I__7921 (
            .O(N__33656),
            .I(N__33646));
    LocalMux I__7920 (
            .O(N__33653),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    LocalMux I__7919 (
            .O(N__33646),
            .I(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ));
    CascadeMux I__7918 (
            .O(N__33641),
            .I(N__33637));
    InMux I__7917 (
            .O(N__33640),
            .I(N__33632));
    InMux I__7916 (
            .O(N__33637),
            .I(N__33625));
    InMux I__7915 (
            .O(N__33636),
            .I(N__33625));
    InMux I__7914 (
            .O(N__33635),
            .I(N__33625));
    LocalMux I__7913 (
            .O(N__33632),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    LocalMux I__7912 (
            .O(N__33625),
            .I(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ));
    CascadeMux I__7911 (
            .O(N__33620),
            .I(N__33617));
    InMux I__7910 (
            .O(N__33617),
            .I(N__33602));
    InMux I__7909 (
            .O(N__33616),
            .I(N__33602));
    InMux I__7908 (
            .O(N__33615),
            .I(N__33599));
    InMux I__7907 (
            .O(N__33614),
            .I(N__33596));
    InMux I__7906 (
            .O(N__33613),
            .I(N__33591));
    InMux I__7905 (
            .O(N__33612),
            .I(N__33588));
    InMux I__7904 (
            .O(N__33611),
            .I(N__33583));
    InMux I__7903 (
            .O(N__33610),
            .I(N__33583));
    InMux I__7902 (
            .O(N__33609),
            .I(N__33579));
    InMux I__7901 (
            .O(N__33608),
            .I(N__33574));
    InMux I__7900 (
            .O(N__33607),
            .I(N__33574));
    LocalMux I__7899 (
            .O(N__33602),
            .I(N__33569));
    LocalMux I__7898 (
            .O(N__33599),
            .I(N__33564));
    LocalMux I__7897 (
            .O(N__33596),
            .I(N__33564));
    InMux I__7896 (
            .O(N__33595),
            .I(N__33561));
    InMux I__7895 (
            .O(N__33594),
            .I(N__33558));
    LocalMux I__7894 (
            .O(N__33591),
            .I(N__33555));
    LocalMux I__7893 (
            .O(N__33588),
            .I(N__33550));
    LocalMux I__7892 (
            .O(N__33583),
            .I(N__33550));
    CascadeMux I__7891 (
            .O(N__33582),
            .I(N__33547));
    LocalMux I__7890 (
            .O(N__33579),
            .I(N__33540));
    LocalMux I__7889 (
            .O(N__33574),
            .I(N__33540));
    CascadeMux I__7888 (
            .O(N__33573),
            .I(N__33537));
    CascadeMux I__7887 (
            .O(N__33572),
            .I(N__33533));
    Span4Mux_h I__7886 (
            .O(N__33569),
            .I(N__33529));
    Span12Mux_v I__7885 (
            .O(N__33564),
            .I(N__33524));
    LocalMux I__7884 (
            .O(N__33561),
            .I(N__33524));
    LocalMux I__7883 (
            .O(N__33558),
            .I(N__33517));
    Span4Mux_v I__7882 (
            .O(N__33555),
            .I(N__33517));
    Span4Mux_h I__7881 (
            .O(N__33550),
            .I(N__33517));
    InMux I__7880 (
            .O(N__33547),
            .I(N__33510));
    InMux I__7879 (
            .O(N__33546),
            .I(N__33510));
    InMux I__7878 (
            .O(N__33545),
            .I(N__33510));
    Span4Mux_h I__7877 (
            .O(N__33540),
            .I(N__33507));
    InMux I__7876 (
            .O(N__33537),
            .I(N__33504));
    InMux I__7875 (
            .O(N__33536),
            .I(N__33499));
    InMux I__7874 (
            .O(N__33533),
            .I(N__33499));
    InMux I__7873 (
            .O(N__33532),
            .I(N__33496));
    Odrv4 I__7872 (
            .O(N__33529),
            .I(\this_vga_signals.vaddress_7 ));
    Odrv12 I__7871 (
            .O(N__33524),
            .I(\this_vga_signals.vaddress_7 ));
    Odrv4 I__7870 (
            .O(N__33517),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__7869 (
            .O(N__33510),
            .I(\this_vga_signals.vaddress_7 ));
    Odrv4 I__7868 (
            .O(N__33507),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__7867 (
            .O(N__33504),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__7866 (
            .O(N__33499),
            .I(\this_vga_signals.vaddress_7 ));
    LocalMux I__7865 (
            .O(N__33496),
            .I(\this_vga_signals.vaddress_7 ));
    InMux I__7864 (
            .O(N__33479),
            .I(N__33467));
    InMux I__7863 (
            .O(N__33478),
            .I(N__33467));
    InMux I__7862 (
            .O(N__33477),
            .I(N__33460));
    InMux I__7861 (
            .O(N__33476),
            .I(N__33460));
    InMux I__7860 (
            .O(N__33475),
            .I(N__33460));
    InMux I__7859 (
            .O(N__33474),
            .I(N__33455));
    InMux I__7858 (
            .O(N__33473),
            .I(N__33455));
    InMux I__7857 (
            .O(N__33472),
            .I(N__33452));
    LocalMux I__7856 (
            .O(N__33467),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__7855 (
            .O(N__33460),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__7854 (
            .O(N__33455),
            .I(\this_vga_signals.vaddress_6 ));
    LocalMux I__7853 (
            .O(N__33452),
            .I(\this_vga_signals.vaddress_6 ));
    InMux I__7852 (
            .O(N__33443),
            .I(N__33436));
    InMux I__7851 (
            .O(N__33442),
            .I(N__33429));
    InMux I__7850 (
            .O(N__33441),
            .I(N__33429));
    InMux I__7849 (
            .O(N__33440),
            .I(N__33429));
    InMux I__7848 (
            .O(N__33439),
            .I(N__33426));
    LocalMux I__7847 (
            .O(N__33436),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__7846 (
            .O(N__33429),
            .I(\this_vga_signals.vaddress_5 ));
    LocalMux I__7845 (
            .O(N__33426),
            .I(\this_vga_signals.vaddress_5 ));
    CascadeMux I__7844 (
            .O(N__33419),
            .I(\this_vga_signals.vaddress_7_cascade_ ));
    InMux I__7843 (
            .O(N__33416),
            .I(N__33404));
    InMux I__7842 (
            .O(N__33415),
            .I(N__33399));
    InMux I__7841 (
            .O(N__33414),
            .I(N__33399));
    InMux I__7840 (
            .O(N__33413),
            .I(N__33396));
    InMux I__7839 (
            .O(N__33412),
            .I(N__33393));
    InMux I__7838 (
            .O(N__33411),
            .I(N__33390));
    InMux I__7837 (
            .O(N__33410),
            .I(N__33385));
    InMux I__7836 (
            .O(N__33409),
            .I(N__33385));
    InMux I__7835 (
            .O(N__33408),
            .I(N__33381));
    InMux I__7834 (
            .O(N__33407),
            .I(N__33377));
    LocalMux I__7833 (
            .O(N__33404),
            .I(N__33374));
    LocalMux I__7832 (
            .O(N__33399),
            .I(N__33371));
    LocalMux I__7831 (
            .O(N__33396),
            .I(N__33367));
    LocalMux I__7830 (
            .O(N__33393),
            .I(N__33360));
    LocalMux I__7829 (
            .O(N__33390),
            .I(N__33360));
    LocalMux I__7828 (
            .O(N__33385),
            .I(N__33360));
    InMux I__7827 (
            .O(N__33384),
            .I(N__33352));
    LocalMux I__7826 (
            .O(N__33381),
            .I(N__33349));
    InMux I__7825 (
            .O(N__33380),
            .I(N__33346));
    LocalMux I__7824 (
            .O(N__33377),
            .I(N__33343));
    Span4Mux_h I__7823 (
            .O(N__33374),
            .I(N__33338));
    Span4Mux_h I__7822 (
            .O(N__33371),
            .I(N__33338));
    InMux I__7821 (
            .O(N__33370),
            .I(N__33335));
    Span4Mux_v I__7820 (
            .O(N__33367),
            .I(N__33330));
    Span4Mux_h I__7819 (
            .O(N__33360),
            .I(N__33330));
    InMux I__7818 (
            .O(N__33359),
            .I(N__33325));
    InMux I__7817 (
            .O(N__33358),
            .I(N__33325));
    InMux I__7816 (
            .O(N__33357),
            .I(N__33320));
    InMux I__7815 (
            .O(N__33356),
            .I(N__33320));
    InMux I__7814 (
            .O(N__33355),
            .I(N__33317));
    LocalMux I__7813 (
            .O(N__33352),
            .I(\this_vga_signals.SUM_2 ));
    Odrv4 I__7812 (
            .O(N__33349),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__7811 (
            .O(N__33346),
            .I(\this_vga_signals.SUM_2 ));
    Odrv4 I__7810 (
            .O(N__33343),
            .I(\this_vga_signals.SUM_2 ));
    Odrv4 I__7809 (
            .O(N__33338),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__7808 (
            .O(N__33335),
            .I(\this_vga_signals.SUM_2 ));
    Odrv4 I__7807 (
            .O(N__33330),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__7806 (
            .O(N__33325),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__7805 (
            .O(N__33320),
            .I(\this_vga_signals.SUM_2 ));
    LocalMux I__7804 (
            .O(N__33317),
            .I(\this_vga_signals.SUM_2 ));
    InMux I__7803 (
            .O(N__33296),
            .I(N__33289));
    InMux I__7802 (
            .O(N__33295),
            .I(N__33284));
    InMux I__7801 (
            .O(N__33294),
            .I(N__33284));
    InMux I__7800 (
            .O(N__33293),
            .I(N__33279));
    InMux I__7799 (
            .O(N__33292),
            .I(N__33279));
    LocalMux I__7798 (
            .O(N__33289),
            .I(\this_vga_signals.if_m2_0 ));
    LocalMux I__7797 (
            .O(N__33284),
            .I(\this_vga_signals.if_m2_0 ));
    LocalMux I__7796 (
            .O(N__33279),
            .I(\this_vga_signals.if_m2_0 ));
    CascadeMux I__7795 (
            .O(N__33272),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_ ));
    CascadeMux I__7794 (
            .O(N__33269),
            .I(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ));
    CascadeMux I__7793 (
            .O(N__33266),
            .I(N__33262));
    InMux I__7792 (
            .O(N__33265),
            .I(N__33258));
    InMux I__7791 (
            .O(N__33262),
            .I(N__33255));
    InMux I__7790 (
            .O(N__33261),
            .I(N__33250));
    LocalMux I__7789 (
            .O(N__33258),
            .I(N__33245));
    LocalMux I__7788 (
            .O(N__33255),
            .I(N__33245));
    CascadeMux I__7787 (
            .O(N__33254),
            .I(N__33242));
    CascadeMux I__7786 (
            .O(N__33253),
            .I(N__33239));
    LocalMux I__7785 (
            .O(N__33250),
            .I(N__33234));
    Span4Mux_v I__7784 (
            .O(N__33245),
            .I(N__33231));
    InMux I__7783 (
            .O(N__33242),
            .I(N__33222));
    InMux I__7782 (
            .O(N__33239),
            .I(N__33222));
    InMux I__7781 (
            .O(N__33238),
            .I(N__33222));
    InMux I__7780 (
            .O(N__33237),
            .I(N__33222));
    Span4Mux_h I__7779 (
            .O(N__33234),
            .I(N__33219));
    Odrv4 I__7778 (
            .O(N__33231),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    LocalMux I__7777 (
            .O(N__33222),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    Odrv4 I__7776 (
            .O(N__33219),
            .I(\this_vga_signals.mult1_un40_sum_c3_0 ));
    CascadeMux I__7775 (
            .O(N__33212),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_ ));
    CascadeMux I__7774 (
            .O(N__33209),
            .I(N__33206));
    InMux I__7773 (
            .O(N__33206),
            .I(N__33203));
    LocalMux I__7772 (
            .O(N__33203),
            .I(N__33200));
    Span4Mux_h I__7771 (
            .O(N__33200),
            .I(N__33197));
    Odrv4 I__7770 (
            .O(N__33197),
            .I(\this_vga_signals.N_14 ));
    InMux I__7769 (
            .O(N__33194),
            .I(N__33188));
    InMux I__7768 (
            .O(N__33193),
            .I(N__33188));
    LocalMux I__7767 (
            .O(N__33188),
            .I(\this_vga_signals.g1_6 ));
    CascadeMux I__7766 (
            .O(N__33185),
            .I(N__33179));
    InMux I__7765 (
            .O(N__33184),
            .I(N__33176));
    CascadeMux I__7764 (
            .O(N__33183),
            .I(N__33173));
    CascadeMux I__7763 (
            .O(N__33182),
            .I(N__33169));
    InMux I__7762 (
            .O(N__33179),
            .I(N__33165));
    LocalMux I__7761 (
            .O(N__33176),
            .I(N__33162));
    InMux I__7760 (
            .O(N__33173),
            .I(N__33159));
    InMux I__7759 (
            .O(N__33172),
            .I(N__33156));
    InMux I__7758 (
            .O(N__33169),
            .I(N__33153));
    CascadeMux I__7757 (
            .O(N__33168),
            .I(N__33150));
    LocalMux I__7756 (
            .O(N__33165),
            .I(N__33146));
    Span4Mux_h I__7755 (
            .O(N__33162),
            .I(N__33141));
    LocalMux I__7754 (
            .O(N__33159),
            .I(N__33141));
    LocalMux I__7753 (
            .O(N__33156),
            .I(N__33138));
    LocalMux I__7752 (
            .O(N__33153),
            .I(N__33135));
    InMux I__7751 (
            .O(N__33150),
            .I(N__33132));
    CascadeMux I__7750 (
            .O(N__33149),
            .I(N__33128));
    Span4Mux_v I__7749 (
            .O(N__33146),
            .I(N__33109));
    Span4Mux_v I__7748 (
            .O(N__33141),
            .I(N__33109));
    Span4Mux_h I__7747 (
            .O(N__33138),
            .I(N__33109));
    Span4Mux_v I__7746 (
            .O(N__33135),
            .I(N__33109));
    LocalMux I__7745 (
            .O(N__33132),
            .I(N__33109));
    CascadeMux I__7744 (
            .O(N__33131),
            .I(N__33106));
    InMux I__7743 (
            .O(N__33128),
            .I(N__33102));
    InMux I__7742 (
            .O(N__33127),
            .I(N__33097));
    InMux I__7741 (
            .O(N__33126),
            .I(N__33097));
    InMux I__7740 (
            .O(N__33125),
            .I(N__33092));
    InMux I__7739 (
            .O(N__33124),
            .I(N__33092));
    InMux I__7738 (
            .O(N__33123),
            .I(N__33089));
    InMux I__7737 (
            .O(N__33122),
            .I(N__33084));
    InMux I__7736 (
            .O(N__33121),
            .I(N__33084));
    CascadeMux I__7735 (
            .O(N__33120),
            .I(N__33080));
    Span4Mux_h I__7734 (
            .O(N__33109),
            .I(N__33074));
    InMux I__7733 (
            .O(N__33106),
            .I(N__33071));
    InMux I__7732 (
            .O(N__33105),
            .I(N__33068));
    LocalMux I__7731 (
            .O(N__33102),
            .I(N__33065));
    LocalMux I__7730 (
            .O(N__33097),
            .I(N__33062));
    LocalMux I__7729 (
            .O(N__33092),
            .I(N__33059));
    LocalMux I__7728 (
            .O(N__33089),
            .I(N__33054));
    LocalMux I__7727 (
            .O(N__33084),
            .I(N__33054));
    InMux I__7726 (
            .O(N__33083),
            .I(N__33051));
    InMux I__7725 (
            .O(N__33080),
            .I(N__33046));
    InMux I__7724 (
            .O(N__33079),
            .I(N__33046));
    InMux I__7723 (
            .O(N__33078),
            .I(N__33041));
    InMux I__7722 (
            .O(N__33077),
            .I(N__33041));
    Span4Mux_h I__7721 (
            .O(N__33074),
            .I(N__33038));
    LocalMux I__7720 (
            .O(N__33071),
            .I(N__33029));
    LocalMux I__7719 (
            .O(N__33068),
            .I(N__33029));
    Span4Mux_h I__7718 (
            .O(N__33065),
            .I(N__33029));
    Span4Mux_h I__7717 (
            .O(N__33062),
            .I(N__33029));
    Span4Mux_v I__7716 (
            .O(N__33059),
            .I(N__33024));
    Span4Mux_h I__7715 (
            .O(N__33054),
            .I(N__33024));
    LocalMux I__7714 (
            .O(N__33051),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__7713 (
            .O(N__33046),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    LocalMux I__7712 (
            .O(N__33041),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__7711 (
            .O(N__33038),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__7710 (
            .O(N__33029),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    Odrv4 I__7709 (
            .O(N__33024),
            .I(\this_vga_signals.M_vcounter_qZ0Z_5 ));
    CascadeMux I__7708 (
            .O(N__33011),
            .I(\this_vga_signals.N_7_1_0_3_cascade_ ));
    InMux I__7707 (
            .O(N__33008),
            .I(N__33005));
    LocalMux I__7706 (
            .O(N__33005),
            .I(\this_vga_signals.G_5_i_o2_0_1 ));
    InMux I__7705 (
            .O(N__33002),
            .I(N__32997));
    InMux I__7704 (
            .O(N__33001),
            .I(N__32993));
    InMux I__7703 (
            .O(N__33000),
            .I(N__32990));
    LocalMux I__7702 (
            .O(N__32997),
            .I(N__32987));
    InMux I__7701 (
            .O(N__32996),
            .I(N__32980));
    LocalMux I__7700 (
            .O(N__32993),
            .I(N__32977));
    LocalMux I__7699 (
            .O(N__32990),
            .I(N__32974));
    Span4Mux_h I__7698 (
            .O(N__32987),
            .I(N__32971));
    InMux I__7697 (
            .O(N__32986),
            .I(N__32964));
    InMux I__7696 (
            .O(N__32985),
            .I(N__32964));
    InMux I__7695 (
            .O(N__32984),
            .I(N__32964));
    InMux I__7694 (
            .O(N__32983),
            .I(N__32961));
    LocalMux I__7693 (
            .O(N__32980),
            .I(\this_vga_signals.vaddress_8 ));
    Odrv4 I__7692 (
            .O(N__32977),
            .I(\this_vga_signals.vaddress_8 ));
    Odrv4 I__7691 (
            .O(N__32974),
            .I(\this_vga_signals.vaddress_8 ));
    Odrv4 I__7690 (
            .O(N__32971),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__7689 (
            .O(N__32964),
            .I(\this_vga_signals.vaddress_8 ));
    LocalMux I__7688 (
            .O(N__32961),
            .I(\this_vga_signals.vaddress_8 ));
    InMux I__7687 (
            .O(N__32948),
            .I(N__32945));
    LocalMux I__7686 (
            .O(N__32945),
            .I(N__32939));
    InMux I__7685 (
            .O(N__32944),
            .I(N__32936));
    CascadeMux I__7684 (
            .O(N__32943),
            .I(N__32931));
    InMux I__7683 (
            .O(N__32942),
            .I(N__32926));
    Span4Mux_v I__7682 (
            .O(N__32939),
            .I(N__32923));
    LocalMux I__7681 (
            .O(N__32936),
            .I(N__32920));
    InMux I__7680 (
            .O(N__32935),
            .I(N__32917));
    InMux I__7679 (
            .O(N__32934),
            .I(N__32914));
    InMux I__7678 (
            .O(N__32931),
            .I(N__32909));
    InMux I__7677 (
            .O(N__32930),
            .I(N__32909));
    InMux I__7676 (
            .O(N__32929),
            .I(N__32906));
    LocalMux I__7675 (
            .O(N__32926),
            .I(\this_vga_signals.vaddress_9 ));
    Odrv4 I__7674 (
            .O(N__32923),
            .I(\this_vga_signals.vaddress_9 ));
    Odrv4 I__7673 (
            .O(N__32920),
            .I(\this_vga_signals.vaddress_9 ));
    LocalMux I__7672 (
            .O(N__32917),
            .I(\this_vga_signals.vaddress_9 ));
    LocalMux I__7671 (
            .O(N__32914),
            .I(\this_vga_signals.vaddress_9 ));
    LocalMux I__7670 (
            .O(N__32909),
            .I(\this_vga_signals.vaddress_9 ));
    LocalMux I__7669 (
            .O(N__32906),
            .I(\this_vga_signals.vaddress_9 ));
    InMux I__7668 (
            .O(N__32891),
            .I(N__32888));
    LocalMux I__7667 (
            .O(N__32888),
            .I(N__32885));
    Odrv4 I__7666 (
            .O(N__32885),
            .I(\this_vga_signals.N_19_0_0 ));
    InMux I__7665 (
            .O(N__32882),
            .I(N__32876));
    InMux I__7664 (
            .O(N__32881),
            .I(N__32873));
    InMux I__7663 (
            .O(N__32880),
            .I(N__32868));
    InMux I__7662 (
            .O(N__32879),
            .I(N__32868));
    LocalMux I__7661 (
            .O(N__32876),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__7660 (
            .O(N__32873),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    LocalMux I__7659 (
            .O(N__32868),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ));
    CascadeMux I__7658 (
            .O(N__32861),
            .I(N__32857));
    CascadeMux I__7657 (
            .O(N__32860),
            .I(N__32851));
    InMux I__7656 (
            .O(N__32857),
            .I(N__32846));
    InMux I__7655 (
            .O(N__32856),
            .I(N__32846));
    InMux I__7654 (
            .O(N__32855),
            .I(N__32843));
    InMux I__7653 (
            .O(N__32854),
            .I(N__32838));
    InMux I__7652 (
            .O(N__32851),
            .I(N__32838));
    LocalMux I__7651 (
            .O(N__32846),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    LocalMux I__7650 (
            .O(N__32843),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    LocalMux I__7649 (
            .O(N__32838),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ));
    InMux I__7648 (
            .O(N__32831),
            .I(N__32827));
    InMux I__7647 (
            .O(N__32830),
            .I(N__32824));
    LocalMux I__7646 (
            .O(N__32827),
            .I(\this_vga_signals.m47_0_0 ));
    LocalMux I__7645 (
            .O(N__32824),
            .I(\this_vga_signals.m47_0_0 ));
    InMux I__7644 (
            .O(N__32819),
            .I(N__32811));
    InMux I__7643 (
            .O(N__32818),
            .I(N__32808));
    InMux I__7642 (
            .O(N__32817),
            .I(N__32805));
    InMux I__7641 (
            .O(N__32816),
            .I(N__32802));
    InMux I__7640 (
            .O(N__32815),
            .I(N__32798));
    InMux I__7639 (
            .O(N__32814),
            .I(N__32795));
    LocalMux I__7638 (
            .O(N__32811),
            .I(N__32790));
    LocalMux I__7637 (
            .O(N__32808),
            .I(N__32790));
    LocalMux I__7636 (
            .O(N__32805),
            .I(N__32785));
    LocalMux I__7635 (
            .O(N__32802),
            .I(N__32785));
    InMux I__7634 (
            .O(N__32801),
            .I(N__32782));
    LocalMux I__7633 (
            .O(N__32798),
            .I(N__32779));
    LocalMux I__7632 (
            .O(N__32795),
            .I(N__32776));
    Span12Mux_s6_v I__7631 (
            .O(N__32790),
            .I(N__32772));
    Span12Mux_v I__7630 (
            .O(N__32785),
            .I(N__32769));
    LocalMux I__7629 (
            .O(N__32782),
            .I(N__32766));
    Span4Mux_h I__7628 (
            .O(N__32779),
            .I(N__32763));
    Span12Mux_h I__7627 (
            .O(N__32776),
            .I(N__32760));
    InMux I__7626 (
            .O(N__32775),
            .I(N__32757));
    Span12Mux_h I__7625 (
            .O(N__32772),
            .I(N__32750));
    Span12Mux_h I__7624 (
            .O(N__32769),
            .I(N__32750));
    Span12Mux_h I__7623 (
            .O(N__32766),
            .I(N__32750));
    Span4Mux_h I__7622 (
            .O(N__32763),
            .I(N__32747));
    Span12Mux_v I__7621 (
            .O(N__32760),
            .I(N__32742));
    LocalMux I__7620 (
            .O(N__32757),
            .I(N__32742));
    Odrv12 I__7619 (
            .O(N__32750),
            .I(M_this_spr_ram_write_data_3));
    Odrv4 I__7618 (
            .O(N__32747),
            .I(M_this_spr_ram_write_data_3));
    Odrv12 I__7617 (
            .O(N__32742),
            .I(M_this_spr_ram_write_data_3));
    InMux I__7616 (
            .O(N__32735),
            .I(N__32732));
    LocalMux I__7615 (
            .O(N__32732),
            .I(N__32729));
    Span4Mux_h I__7614 (
            .O(N__32729),
            .I(N__32726));
    Odrv4 I__7613 (
            .O(N__32726),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_1 ));
    InMux I__7612 (
            .O(N__32723),
            .I(N__32720));
    LocalMux I__7611 (
            .O(N__32720),
            .I(N__32717));
    Span4Mux_v I__7610 (
            .O(N__32717),
            .I(N__32714));
    Span4Mux_v I__7609 (
            .O(N__32714),
            .I(N__32711));
    Span4Mux_h I__7608 (
            .O(N__32711),
            .I(N__32708));
    Odrv4 I__7607 (
            .O(N__32708),
            .I(M_this_map_ram_read_data_1));
    CascadeMux I__7606 (
            .O(N__32705),
            .I(N__32702));
    InMux I__7605 (
            .O(N__32702),
            .I(N__32698));
    InMux I__7604 (
            .O(N__32701),
            .I(N__32695));
    LocalMux I__7603 (
            .O(N__32698),
            .I(N__32690));
    LocalMux I__7602 (
            .O(N__32695),
            .I(N__32684));
    InMux I__7601 (
            .O(N__32694),
            .I(N__32681));
    InMux I__7600 (
            .O(N__32693),
            .I(N__32677));
    Span4Mux_h I__7599 (
            .O(N__32690),
            .I(N__32674));
    InMux I__7598 (
            .O(N__32689),
            .I(N__32671));
    InMux I__7597 (
            .O(N__32688),
            .I(N__32666));
    InMux I__7596 (
            .O(N__32687),
            .I(N__32660));
    Span4Mux_h I__7595 (
            .O(N__32684),
            .I(N__32655));
    LocalMux I__7594 (
            .O(N__32681),
            .I(N__32655));
    InMux I__7593 (
            .O(N__32680),
            .I(N__32652));
    LocalMux I__7592 (
            .O(N__32677),
            .I(N__32649));
    Span4Mux_h I__7591 (
            .O(N__32674),
            .I(N__32644));
    LocalMux I__7590 (
            .O(N__32671),
            .I(N__32644));
    InMux I__7589 (
            .O(N__32670),
            .I(N__32641));
    InMux I__7588 (
            .O(N__32669),
            .I(N__32638));
    LocalMux I__7587 (
            .O(N__32666),
            .I(N__32635));
    InMux I__7586 (
            .O(N__32665),
            .I(N__32632));
    InMux I__7585 (
            .O(N__32664),
            .I(N__32627));
    InMux I__7584 (
            .O(N__32663),
            .I(N__32627));
    LocalMux I__7583 (
            .O(N__32660),
            .I(N__32620));
    Span4Mux_v I__7582 (
            .O(N__32655),
            .I(N__32620));
    LocalMux I__7581 (
            .O(N__32652),
            .I(N__32620));
    Span4Mux_v I__7580 (
            .O(N__32649),
            .I(N__32617));
    Sp12to4 I__7579 (
            .O(N__32644),
            .I(N__32612));
    LocalMux I__7578 (
            .O(N__32641),
            .I(N__32612));
    LocalMux I__7577 (
            .O(N__32638),
            .I(N__32603));
    Span4Mux_h I__7576 (
            .O(N__32635),
            .I(N__32603));
    LocalMux I__7575 (
            .O(N__32632),
            .I(N__32603));
    LocalMux I__7574 (
            .O(N__32627),
            .I(N__32603));
    Span4Mux_h I__7573 (
            .O(N__32620),
            .I(N__32600));
    Sp12to4 I__7572 (
            .O(N__32617),
            .I(N__32595));
    Span12Mux_v I__7571 (
            .O(N__32612),
            .I(N__32595));
    Odrv4 I__7570 (
            .O(N__32603),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv4 I__7569 (
            .O(N__32600),
            .I(\this_ppu.M_state_q_inv_1 ));
    Odrv12 I__7568 (
            .O(N__32595),
            .I(\this_ppu.M_state_q_inv_1 ));
    CascadeMux I__7567 (
            .O(N__32588),
            .I(N__32584));
    CascadeMux I__7566 (
            .O(N__32587),
            .I(N__32581));
    InMux I__7565 (
            .O(N__32584),
            .I(N__32575));
    InMux I__7564 (
            .O(N__32581),
            .I(N__32572));
    CascadeMux I__7563 (
            .O(N__32580),
            .I(N__32569));
    CascadeMux I__7562 (
            .O(N__32579),
            .I(N__32566));
    CascadeMux I__7561 (
            .O(N__32578),
            .I(N__32558));
    LocalMux I__7560 (
            .O(N__32575),
            .I(N__32550));
    LocalMux I__7559 (
            .O(N__32572),
            .I(N__32550));
    InMux I__7558 (
            .O(N__32569),
            .I(N__32547));
    InMux I__7557 (
            .O(N__32566),
            .I(N__32544));
    CascadeMux I__7556 (
            .O(N__32565),
            .I(N__32541));
    CascadeMux I__7555 (
            .O(N__32564),
            .I(N__32538));
    CascadeMux I__7554 (
            .O(N__32563),
            .I(N__32532));
    CascadeMux I__7553 (
            .O(N__32562),
            .I(N__32529));
    CascadeMux I__7552 (
            .O(N__32561),
            .I(N__32526));
    InMux I__7551 (
            .O(N__32558),
            .I(N__32523));
    CascadeMux I__7550 (
            .O(N__32557),
            .I(N__32520));
    CascadeMux I__7549 (
            .O(N__32556),
            .I(N__32517));
    CascadeMux I__7548 (
            .O(N__32555),
            .I(N__32514));
    Span4Mux_s3_v I__7547 (
            .O(N__32550),
            .I(N__32507));
    LocalMux I__7546 (
            .O(N__32547),
            .I(N__32507));
    LocalMux I__7545 (
            .O(N__32544),
            .I(N__32507));
    InMux I__7544 (
            .O(N__32541),
            .I(N__32504));
    InMux I__7543 (
            .O(N__32538),
            .I(N__32501));
    CascadeMux I__7542 (
            .O(N__32537),
            .I(N__32498));
    CascadeMux I__7541 (
            .O(N__32536),
            .I(N__32495));
    CascadeMux I__7540 (
            .O(N__32535),
            .I(N__32492));
    InMux I__7539 (
            .O(N__32532),
            .I(N__32489));
    InMux I__7538 (
            .O(N__32529),
            .I(N__32486));
    InMux I__7537 (
            .O(N__32526),
            .I(N__32483));
    LocalMux I__7536 (
            .O(N__32523),
            .I(N__32480));
    InMux I__7535 (
            .O(N__32520),
            .I(N__32477));
    InMux I__7534 (
            .O(N__32517),
            .I(N__32474));
    InMux I__7533 (
            .O(N__32514),
            .I(N__32471));
    Span4Mux_v I__7532 (
            .O(N__32507),
            .I(N__32464));
    LocalMux I__7531 (
            .O(N__32504),
            .I(N__32464));
    LocalMux I__7530 (
            .O(N__32501),
            .I(N__32464));
    InMux I__7529 (
            .O(N__32498),
            .I(N__32461));
    InMux I__7528 (
            .O(N__32495),
            .I(N__32458));
    InMux I__7527 (
            .O(N__32492),
            .I(N__32455));
    LocalMux I__7526 (
            .O(N__32489),
            .I(N__32452));
    LocalMux I__7525 (
            .O(N__32486),
            .I(N__32447));
    LocalMux I__7524 (
            .O(N__32483),
            .I(N__32447));
    Span12Mux_s7_v I__7523 (
            .O(N__32480),
            .I(N__32440));
    LocalMux I__7522 (
            .O(N__32477),
            .I(N__32440));
    LocalMux I__7521 (
            .O(N__32474),
            .I(N__32440));
    LocalMux I__7520 (
            .O(N__32471),
            .I(N__32437));
    Span4Mux_v I__7519 (
            .O(N__32464),
            .I(N__32430));
    LocalMux I__7518 (
            .O(N__32461),
            .I(N__32430));
    LocalMux I__7517 (
            .O(N__32458),
            .I(N__32430));
    LocalMux I__7516 (
            .O(N__32455),
            .I(N__32427));
    Span12Mux_h I__7515 (
            .O(N__32452),
            .I(N__32424));
    Span12Mux_v I__7514 (
            .O(N__32447),
            .I(N__32419));
    Span12Mux_v I__7513 (
            .O(N__32440),
            .I(N__32419));
    Span4Mux_v I__7512 (
            .O(N__32437),
            .I(N__32414));
    Span4Mux_v I__7511 (
            .O(N__32430),
            .I(N__32414));
    Span12Mux_h I__7510 (
            .O(N__32427),
            .I(N__32411));
    Span12Mux_v I__7509 (
            .O(N__32424),
            .I(N__32406));
    Span12Mux_h I__7508 (
            .O(N__32419),
            .I(N__32406));
    Span4Mux_h I__7507 (
            .O(N__32414),
            .I(N__32403));
    Odrv12 I__7506 (
            .O(N__32411),
            .I(M_this_ppu_spr_addr_7));
    Odrv12 I__7505 (
            .O(N__32406),
            .I(M_this_ppu_spr_addr_7));
    Odrv4 I__7504 (
            .O(N__32403),
            .I(M_this_ppu_spr_addr_7));
    InMux I__7503 (
            .O(N__32396),
            .I(N__32393));
    LocalMux I__7502 (
            .O(N__32393),
            .I(N__32389));
    InMux I__7501 (
            .O(N__32392),
            .I(N__32386));
    Span4Mux_h I__7500 (
            .O(N__32389),
            .I(N__32382));
    LocalMux I__7499 (
            .O(N__32386),
            .I(N__32379));
    InMux I__7498 (
            .O(N__32385),
            .I(N__32376));
    Span4Mux_v I__7497 (
            .O(N__32382),
            .I(N__32367));
    Span4Mux_h I__7496 (
            .O(N__32379),
            .I(N__32367));
    LocalMux I__7495 (
            .O(N__32376),
            .I(N__32364));
    InMux I__7494 (
            .O(N__32375),
            .I(N__32361));
    InMux I__7493 (
            .O(N__32374),
            .I(N__32357));
    InMux I__7492 (
            .O(N__32373),
            .I(N__32354));
    InMux I__7491 (
            .O(N__32372),
            .I(N__32351));
    Span4Mux_v I__7490 (
            .O(N__32367),
            .I(N__32346));
    Span4Mux_h I__7489 (
            .O(N__32364),
            .I(N__32346));
    LocalMux I__7488 (
            .O(N__32361),
            .I(N__32343));
    InMux I__7487 (
            .O(N__32360),
            .I(N__32340));
    LocalMux I__7486 (
            .O(N__32357),
            .I(N__32335));
    LocalMux I__7485 (
            .O(N__32354),
            .I(N__32335));
    LocalMux I__7484 (
            .O(N__32351),
            .I(N__32332));
    Span4Mux_v I__7483 (
            .O(N__32346),
            .I(N__32327));
    Span4Mux_h I__7482 (
            .O(N__32343),
            .I(N__32327));
    LocalMux I__7481 (
            .O(N__32340),
            .I(N__32324));
    Span12Mux_s10_v I__7480 (
            .O(N__32335),
            .I(N__32321));
    Span12Mux_s9_v I__7479 (
            .O(N__32332),
            .I(N__32318));
    Span4Mux_v I__7478 (
            .O(N__32327),
            .I(N__32313));
    Span4Mux_h I__7477 (
            .O(N__32324),
            .I(N__32313));
    Span12Mux_h I__7476 (
            .O(N__32321),
            .I(N__32308));
    Span12Mux_h I__7475 (
            .O(N__32318),
            .I(N__32308));
    Span4Mux_h I__7474 (
            .O(N__32313),
            .I(N__32305));
    Odrv12 I__7473 (
            .O(N__32308),
            .I(M_this_spr_ram_write_data_1));
    Odrv4 I__7472 (
            .O(N__32305),
            .I(M_this_spr_ram_write_data_1));
    CascadeMux I__7471 (
            .O(N__32300),
            .I(M_this_state_d_0_sqmuxa_2_cascade_));
    CascadeMux I__7470 (
            .O(N__32297),
            .I(\this_start_data_delay.N_233_0_cascade_ ));
    CEMux I__7469 (
            .O(N__32294),
            .I(N__32291));
    LocalMux I__7468 (
            .O(N__32291),
            .I(N__32287));
    CEMux I__7467 (
            .O(N__32290),
            .I(N__32283));
    Span4Mux_h I__7466 (
            .O(N__32287),
            .I(N__32280));
    CEMux I__7465 (
            .O(N__32286),
            .I(N__32277));
    LocalMux I__7464 (
            .O(N__32283),
            .I(N__32270));
    Span4Mux_h I__7463 (
            .O(N__32280),
            .I(N__32270));
    LocalMux I__7462 (
            .O(N__32277),
            .I(N__32270));
    Span4Mux_h I__7461 (
            .O(N__32270),
            .I(N__32267));
    Odrv4 I__7460 (
            .O(N__32267),
            .I(N_164));
    InMux I__7459 (
            .O(N__32264),
            .I(N__32261));
    LocalMux I__7458 (
            .O(N__32261),
            .I(N__32258));
    Span4Mux_v I__7457 (
            .O(N__32258),
            .I(N__32255));
    Odrv4 I__7456 (
            .O(N__32255),
            .I(\this_vga_signals.g1_3_0 ));
    InMux I__7455 (
            .O(N__32252),
            .I(N__32249));
    LocalMux I__7454 (
            .O(N__32249),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6 ));
    CEMux I__7453 (
            .O(N__32246),
            .I(N__32242));
    CEMux I__7452 (
            .O(N__32245),
            .I(N__32239));
    LocalMux I__7451 (
            .O(N__32242),
            .I(N__32236));
    LocalMux I__7450 (
            .O(N__32239),
            .I(N__32233));
    Span4Mux_v I__7449 (
            .O(N__32236),
            .I(N__32228));
    Span4Mux_v I__7448 (
            .O(N__32233),
            .I(N__32228));
    Span4Mux_h I__7447 (
            .O(N__32228),
            .I(N__32225));
    Odrv4 I__7446 (
            .O(N__32225),
            .I(\this_spr_ram.mem_WE_6 ));
    InMux I__7445 (
            .O(N__32222),
            .I(N__32219));
    LocalMux I__7444 (
            .O(N__32219),
            .I(N__32214));
    InMux I__7443 (
            .O(N__32218),
            .I(N__32210));
    InMux I__7442 (
            .O(N__32217),
            .I(N__32206));
    Span4Mux_v I__7441 (
            .O(N__32214),
            .I(N__32201));
    InMux I__7440 (
            .O(N__32213),
            .I(N__32198));
    LocalMux I__7439 (
            .O(N__32210),
            .I(N__32195));
    InMux I__7438 (
            .O(N__32209),
            .I(N__32192));
    LocalMux I__7437 (
            .O(N__32206),
            .I(N__32189));
    InMux I__7436 (
            .O(N__32205),
            .I(N__32186));
    InMux I__7435 (
            .O(N__32204),
            .I(N__32183));
    Span4Mux_v I__7434 (
            .O(N__32201),
            .I(N__32178));
    LocalMux I__7433 (
            .O(N__32198),
            .I(N__32178));
    Span4Mux_h I__7432 (
            .O(N__32195),
            .I(N__32173));
    LocalMux I__7431 (
            .O(N__32192),
            .I(N__32170));
    Span4Mux_h I__7430 (
            .O(N__32189),
            .I(N__32167));
    LocalMux I__7429 (
            .O(N__32186),
            .I(N__32164));
    LocalMux I__7428 (
            .O(N__32183),
            .I(N__32161));
    Span4Mux_v I__7427 (
            .O(N__32178),
            .I(N__32158));
    InMux I__7426 (
            .O(N__32177),
            .I(N__32155));
    InMux I__7425 (
            .O(N__32176),
            .I(N__32152));
    Span4Mux_h I__7424 (
            .O(N__32173),
            .I(N__32147));
    Span4Mux_v I__7423 (
            .O(N__32170),
            .I(N__32147));
    Span4Mux_v I__7422 (
            .O(N__32167),
            .I(N__32140));
    Span4Mux_h I__7421 (
            .O(N__32164),
            .I(N__32140));
    Span4Mux_h I__7420 (
            .O(N__32161),
            .I(N__32140));
    Sp12to4 I__7419 (
            .O(N__32158),
            .I(N__32135));
    LocalMux I__7418 (
            .O(N__32155),
            .I(N__32135));
    LocalMux I__7417 (
            .O(N__32152),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__7416 (
            .O(N__32147),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv4 I__7415 (
            .O(N__32140),
            .I(M_this_spr_address_qZ0Z_12));
    Odrv12 I__7414 (
            .O(N__32135),
            .I(M_this_spr_address_qZ0Z_12));
    InMux I__7413 (
            .O(N__32126),
            .I(N__32122));
    InMux I__7412 (
            .O(N__32125),
            .I(N__32119));
    LocalMux I__7411 (
            .O(N__32122),
            .I(N__32113));
    LocalMux I__7410 (
            .O(N__32119),
            .I(N__32110));
    InMux I__7409 (
            .O(N__32118),
            .I(N__32107));
    InMux I__7408 (
            .O(N__32117),
            .I(N__32104));
    InMux I__7407 (
            .O(N__32116),
            .I(N__32099));
    Span4Mux_v I__7406 (
            .O(N__32113),
            .I(N__32094));
    Span4Mux_h I__7405 (
            .O(N__32110),
            .I(N__32094));
    LocalMux I__7404 (
            .O(N__32107),
            .I(N__32091));
    LocalMux I__7403 (
            .O(N__32104),
            .I(N__32088));
    InMux I__7402 (
            .O(N__32103),
            .I(N__32085));
    InMux I__7401 (
            .O(N__32102),
            .I(N__32082));
    LocalMux I__7400 (
            .O(N__32099),
            .I(N__32077));
    Span4Mux_v I__7399 (
            .O(N__32094),
            .I(N__32072));
    Span4Mux_v I__7398 (
            .O(N__32091),
            .I(N__32072));
    Span4Mux_v I__7397 (
            .O(N__32088),
            .I(N__32067));
    LocalMux I__7396 (
            .O(N__32085),
            .I(N__32067));
    LocalMux I__7395 (
            .O(N__32082),
            .I(N__32064));
    InMux I__7394 (
            .O(N__32081),
            .I(N__32061));
    InMux I__7393 (
            .O(N__32080),
            .I(N__32058));
    Span4Mux_v I__7392 (
            .O(N__32077),
            .I(N__32055));
    Span4Mux_h I__7391 (
            .O(N__32072),
            .I(N__32048));
    Span4Mux_v I__7390 (
            .O(N__32067),
            .I(N__32048));
    Span4Mux_v I__7389 (
            .O(N__32064),
            .I(N__32048));
    LocalMux I__7388 (
            .O(N__32061),
            .I(N__32045));
    LocalMux I__7387 (
            .O(N__32058),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__7386 (
            .O(N__32055),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__7385 (
            .O(N__32048),
            .I(M_this_spr_address_qZ0Z_11));
    Odrv4 I__7384 (
            .O(N__32045),
            .I(M_this_spr_address_qZ0Z_11));
    CascadeMux I__7383 (
            .O(N__32036),
            .I(N__32033));
    InMux I__7382 (
            .O(N__32033),
            .I(N__32027));
    CascadeMux I__7381 (
            .O(N__32032),
            .I(N__32024));
    CascadeMux I__7380 (
            .O(N__32031),
            .I(N__32021));
    CascadeMux I__7379 (
            .O(N__32030),
            .I(N__32018));
    LocalMux I__7378 (
            .O(N__32027),
            .I(N__32013));
    InMux I__7377 (
            .O(N__32024),
            .I(N__32010));
    InMux I__7376 (
            .O(N__32021),
            .I(N__32007));
    InMux I__7375 (
            .O(N__32018),
            .I(N__32004));
    CascadeMux I__7374 (
            .O(N__32017),
            .I(N__32001));
    CascadeMux I__7373 (
            .O(N__32016),
            .I(N__31997));
    Span4Mux_v I__7372 (
            .O(N__32013),
            .I(N__31991));
    LocalMux I__7371 (
            .O(N__32010),
            .I(N__31991));
    LocalMux I__7370 (
            .O(N__32007),
            .I(N__31988));
    LocalMux I__7369 (
            .O(N__32004),
            .I(N__31985));
    InMux I__7368 (
            .O(N__32001),
            .I(N__31982));
    InMux I__7367 (
            .O(N__32000),
            .I(N__31979));
    InMux I__7366 (
            .O(N__31997),
            .I(N__31976));
    CascadeMux I__7365 (
            .O(N__31996),
            .I(N__31973));
    Span4Mux_h I__7364 (
            .O(N__31991),
            .I(N__31969));
    Span4Mux_v I__7363 (
            .O(N__31988),
            .I(N__31966));
    Span4Mux_v I__7362 (
            .O(N__31985),
            .I(N__31963));
    LocalMux I__7361 (
            .O(N__31982),
            .I(N__31960));
    LocalMux I__7360 (
            .O(N__31979),
            .I(N__31957));
    LocalMux I__7359 (
            .O(N__31976),
            .I(N__31954));
    InMux I__7358 (
            .O(N__31973),
            .I(N__31951));
    InMux I__7357 (
            .O(N__31972),
            .I(N__31948));
    Span4Mux_v I__7356 (
            .O(N__31969),
            .I(N__31941));
    Span4Mux_v I__7355 (
            .O(N__31966),
            .I(N__31941));
    Span4Mux_h I__7354 (
            .O(N__31963),
            .I(N__31941));
    Span4Mux_v I__7353 (
            .O(N__31960),
            .I(N__31938));
    Span4Mux_h I__7352 (
            .O(N__31957),
            .I(N__31935));
    Span4Mux_v I__7351 (
            .O(N__31954),
            .I(N__31930));
    LocalMux I__7350 (
            .O(N__31951),
            .I(N__31930));
    LocalMux I__7349 (
            .O(N__31948),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__7348 (
            .O(N__31941),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__7347 (
            .O(N__31938),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__7346 (
            .O(N__31935),
            .I(M_this_spr_address_qZ0Z_13));
    Odrv4 I__7345 (
            .O(N__31930),
            .I(M_this_spr_address_qZ0Z_13));
    InMux I__7344 (
            .O(N__31919),
            .I(N__31915));
    InMux I__7343 (
            .O(N__31918),
            .I(N__31908));
    LocalMux I__7342 (
            .O(N__31915),
            .I(N__31905));
    InMux I__7341 (
            .O(N__31914),
            .I(N__31902));
    InMux I__7340 (
            .O(N__31913),
            .I(N__31899));
    InMux I__7339 (
            .O(N__31912),
            .I(N__31895));
    InMux I__7338 (
            .O(N__31911),
            .I(N__31892));
    LocalMux I__7337 (
            .O(N__31908),
            .I(N__31889));
    Span4Mux_v I__7336 (
            .O(N__31905),
            .I(N__31884));
    LocalMux I__7335 (
            .O(N__31902),
            .I(N__31884));
    LocalMux I__7334 (
            .O(N__31899),
            .I(N__31881));
    InMux I__7333 (
            .O(N__31898),
            .I(N__31878));
    LocalMux I__7332 (
            .O(N__31895),
            .I(N__31873));
    LocalMux I__7331 (
            .O(N__31892),
            .I(N__31873));
    Span4Mux_h I__7330 (
            .O(N__31889),
            .I(N__31870));
    Span4Mux_h I__7329 (
            .O(N__31884),
            .I(N__31867));
    Span4Mux_h I__7328 (
            .O(N__31881),
            .I(N__31864));
    LocalMux I__7327 (
            .O(N__31878),
            .I(N__31861));
    Span12Mux_h I__7326 (
            .O(N__31873),
            .I(N__31858));
    Span4Mux_h I__7325 (
            .O(N__31870),
            .I(N__31855));
    Span4Mux_v I__7324 (
            .O(N__31867),
            .I(N__31850));
    Span4Mux_h I__7323 (
            .O(N__31864),
            .I(N__31850));
    Span4Mux_h I__7322 (
            .O(N__31861),
            .I(N__31847));
    Odrv12 I__7321 (
            .O(N__31858),
            .I(M_this_spr_ram_write_en_0_i_1_0));
    Odrv4 I__7320 (
            .O(N__31855),
            .I(M_this_spr_ram_write_en_0_i_1_0));
    Odrv4 I__7319 (
            .O(N__31850),
            .I(M_this_spr_ram_write_en_0_i_1_0));
    Odrv4 I__7318 (
            .O(N__31847),
            .I(M_this_spr_ram_write_en_0_i_1_0));
    CEMux I__7317 (
            .O(N__31838),
            .I(N__31834));
    CEMux I__7316 (
            .O(N__31837),
            .I(N__31831));
    LocalMux I__7315 (
            .O(N__31834),
            .I(N__31828));
    LocalMux I__7314 (
            .O(N__31831),
            .I(N__31825));
    Span4Mux_v I__7313 (
            .O(N__31828),
            .I(N__31822));
    Span4Mux_h I__7312 (
            .O(N__31825),
            .I(N__31819));
    Span4Mux_h I__7311 (
            .O(N__31822),
            .I(N__31816));
    Span4Mux_h I__7310 (
            .O(N__31819),
            .I(N__31813));
    Odrv4 I__7309 (
            .O(N__31816),
            .I(\this_spr_ram.mem_WE_4 ));
    Odrv4 I__7308 (
            .O(N__31813),
            .I(\this_spr_ram.mem_WE_4 ));
    CascadeMux I__7307 (
            .O(N__31808),
            .I(N__31804));
    InMux I__7306 (
            .O(N__31807),
            .I(N__31801));
    InMux I__7305 (
            .O(N__31804),
            .I(N__31798));
    LocalMux I__7304 (
            .O(N__31801),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ));
    LocalMux I__7303 (
            .O(N__31798),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ));
    InMux I__7302 (
            .O(N__31793),
            .I(N__31790));
    LocalMux I__7301 (
            .O(N__31790),
            .I(\this_vga_signals.mult1_un61_sum_axb1_0_1 ));
    InMux I__7300 (
            .O(N__31787),
            .I(N__31784));
    LocalMux I__7299 (
            .O(N__31784),
            .I(N__31778));
    InMux I__7298 (
            .O(N__31783),
            .I(N__31771));
    InMux I__7297 (
            .O(N__31782),
            .I(N__31771));
    InMux I__7296 (
            .O(N__31781),
            .I(N__31771));
    Odrv4 I__7295 (
            .O(N__31778),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6 ));
    LocalMux I__7294 (
            .O(N__31771),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6 ));
    CascadeMux I__7293 (
            .O(N__31766),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_ ));
    InMux I__7292 (
            .O(N__31763),
            .I(N__31760));
    LocalMux I__7291 (
            .O(N__31760),
            .I(N__31757));
    Odrv4 I__7290 (
            .O(N__31757),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_x0 ));
    InMux I__7289 (
            .O(N__31754),
            .I(N__31746));
    InMux I__7288 (
            .O(N__31753),
            .I(N__31746));
    InMux I__7287 (
            .O(N__31752),
            .I(N__31743));
    InMux I__7286 (
            .O(N__31751),
            .I(N__31740));
    LocalMux I__7285 (
            .O(N__31746),
            .I(N__31732));
    LocalMux I__7284 (
            .O(N__31743),
            .I(N__31727));
    LocalMux I__7283 (
            .O(N__31740),
            .I(N__31727));
    InMux I__7282 (
            .O(N__31739),
            .I(N__31722));
    InMux I__7281 (
            .O(N__31738),
            .I(N__31722));
    InMux I__7280 (
            .O(N__31737),
            .I(N__31711));
    InMux I__7279 (
            .O(N__31736),
            .I(N__31711));
    InMux I__7278 (
            .O(N__31735),
            .I(N__31711));
    Span4Mux_h I__7277 (
            .O(N__31732),
            .I(N__31706));
    Span4Mux_v I__7276 (
            .O(N__31727),
            .I(N__31706));
    LocalMux I__7275 (
            .O(N__31722),
            .I(N__31703));
    InMux I__7274 (
            .O(N__31721),
            .I(N__31700));
    InMux I__7273 (
            .O(N__31720),
            .I(N__31693));
    InMux I__7272 (
            .O(N__31719),
            .I(N__31693));
    InMux I__7271 (
            .O(N__31718),
            .I(N__31693));
    LocalMux I__7270 (
            .O(N__31711),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns ));
    Odrv4 I__7269 (
            .O(N__31706),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns ));
    Odrv12 I__7268 (
            .O(N__31703),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns ));
    LocalMux I__7267 (
            .O(N__31700),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns ));
    LocalMux I__7266 (
            .O(N__31693),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns ));
    CascadeMux I__7265 (
            .O(N__31682),
            .I(\this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_ ));
    InMux I__7264 (
            .O(N__31679),
            .I(N__31672));
    InMux I__7263 (
            .O(N__31678),
            .I(N__31668));
    InMux I__7262 (
            .O(N__31677),
            .I(N__31655));
    InMux I__7261 (
            .O(N__31676),
            .I(N__31655));
    InMux I__7260 (
            .O(N__31675),
            .I(N__31652));
    LocalMux I__7259 (
            .O(N__31672),
            .I(N__31649));
    InMux I__7258 (
            .O(N__31671),
            .I(N__31646));
    LocalMux I__7257 (
            .O(N__31668),
            .I(N__31643));
    InMux I__7256 (
            .O(N__31667),
            .I(N__31640));
    InMux I__7255 (
            .O(N__31666),
            .I(N__31631));
    InMux I__7254 (
            .O(N__31665),
            .I(N__31631));
    InMux I__7253 (
            .O(N__31664),
            .I(N__31631));
    InMux I__7252 (
            .O(N__31663),
            .I(N__31631));
    InMux I__7251 (
            .O(N__31662),
            .I(N__31624));
    InMux I__7250 (
            .O(N__31661),
            .I(N__31624));
    InMux I__7249 (
            .O(N__31660),
            .I(N__31624));
    LocalMux I__7248 (
            .O(N__31655),
            .I(N__31619));
    LocalMux I__7247 (
            .O(N__31652),
            .I(N__31619));
    Odrv4 I__7246 (
            .O(N__31649),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__7245 (
            .O(N__31646),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__7244 (
            .O(N__31643),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__7243 (
            .O(N__31640),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__7242 (
            .O(N__31631),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    LocalMux I__7241 (
            .O(N__31624),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    Odrv4 I__7240 (
            .O(N__31619),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1 ));
    InMux I__7239 (
            .O(N__31604),
            .I(N__31601));
    LocalMux I__7238 (
            .O(N__31601),
            .I(\this_vga_signals.g0_2_0_1 ));
    CascadeMux I__7237 (
            .O(N__31598),
            .I(N__31595));
    InMux I__7236 (
            .O(N__31595),
            .I(N__31588));
    InMux I__7235 (
            .O(N__31594),
            .I(N__31588));
    InMux I__7234 (
            .O(N__31593),
            .I(N__31585));
    LocalMux I__7233 (
            .O(N__31588),
            .I(N__31582));
    LocalMux I__7232 (
            .O(N__31585),
            .I(\this_vga_signals.mult1_un54_sum_axb1_out_0 ));
    Odrv4 I__7231 (
            .O(N__31582),
            .I(\this_vga_signals.mult1_un54_sum_axb1_out_0 ));
    InMux I__7230 (
            .O(N__31577),
            .I(N__31574));
    LocalMux I__7229 (
            .O(N__31574),
            .I(N__31569));
    InMux I__7228 (
            .O(N__31573),
            .I(N__31566));
    InMux I__7227 (
            .O(N__31572),
            .I(N__31563));
    Span4Mux_v I__7226 (
            .O(N__31569),
            .I(N__31556));
    LocalMux I__7225 (
            .O(N__31566),
            .I(N__31556));
    LocalMux I__7224 (
            .O(N__31563),
            .I(N__31556));
    Span4Mux_v I__7223 (
            .O(N__31556),
            .I(N__31553));
    Odrv4 I__7222 (
            .O(N__31553),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ));
    InMux I__7221 (
            .O(N__31550),
            .I(N__31547));
    LocalMux I__7220 (
            .O(N__31547),
            .I(N__31544));
    Sp12to4 I__7219 (
            .O(N__31544),
            .I(N__31541));
    Span12Mux_h I__7218 (
            .O(N__31541),
            .I(N__31537));
    InMux I__7217 (
            .O(N__31540),
            .I(N__31534));
    Odrv12 I__7216 (
            .O(N__31537),
            .I(port_rw_in));
    LocalMux I__7215 (
            .O(N__31534),
            .I(port_rw_in));
    InMux I__7214 (
            .O(N__31529),
            .I(N__31519));
    InMux I__7213 (
            .O(N__31528),
            .I(N__31514));
    InMux I__7212 (
            .O(N__31527),
            .I(N__31514));
    InMux I__7211 (
            .O(N__31526),
            .I(N__31511));
    InMux I__7210 (
            .O(N__31525),
            .I(N__31506));
    InMux I__7209 (
            .O(N__31524),
            .I(N__31506));
    InMux I__7208 (
            .O(N__31523),
            .I(N__31503));
    InMux I__7207 (
            .O(N__31522),
            .I(N__31500));
    LocalMux I__7206 (
            .O(N__31519),
            .I(N__31489));
    LocalMux I__7205 (
            .O(N__31514),
            .I(N__31489));
    LocalMux I__7204 (
            .O(N__31511),
            .I(N__31489));
    LocalMux I__7203 (
            .O(N__31506),
            .I(N__31486));
    LocalMux I__7202 (
            .O(N__31503),
            .I(N__31483));
    LocalMux I__7201 (
            .O(N__31500),
            .I(N__31480));
    InMux I__7200 (
            .O(N__31499),
            .I(N__31477));
    InMux I__7199 (
            .O(N__31498),
            .I(N__31472));
    InMux I__7198 (
            .O(N__31497),
            .I(N__31472));
    InMux I__7197 (
            .O(N__31496),
            .I(N__31469));
    Span4Mux_v I__7196 (
            .O(N__31489),
            .I(N__31466));
    Odrv4 I__7195 (
            .O(N__31486),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__7194 (
            .O(N__31483),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__7193 (
            .O(N__31480),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__7192 (
            .O(N__31477),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__7191 (
            .O(N__31472),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    LocalMux I__7190 (
            .O(N__31469),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    Odrv4 I__7189 (
            .O(N__31466),
            .I(\this_vga_signals.mult1_un47_sum_axbxc1 ));
    InMux I__7188 (
            .O(N__31451),
            .I(N__31448));
    LocalMux I__7187 (
            .O(N__31448),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9 ));
    InMux I__7186 (
            .O(N__31445),
            .I(N__31442));
    LocalMux I__7185 (
            .O(N__31442),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6 ));
    CascadeMux I__7184 (
            .O(N__31439),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_ ));
    CascadeMux I__7183 (
            .O(N__31436),
            .I(\this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_ ));
    InMux I__7182 (
            .O(N__31433),
            .I(N__31430));
    LocalMux I__7181 (
            .O(N__31430),
            .I(\this_vga_signals.g0_5_5 ));
    CascadeMux I__7180 (
            .O(N__31427),
            .I(N__31423));
    InMux I__7179 (
            .O(N__31426),
            .I(N__31416));
    InMux I__7178 (
            .O(N__31423),
            .I(N__31416));
    CascadeMux I__7177 (
            .O(N__31422),
            .I(N__31413));
    CascadeMux I__7176 (
            .O(N__31421),
            .I(N__31402));
    LocalMux I__7175 (
            .O(N__31416),
            .I(N__31396));
    InMux I__7174 (
            .O(N__31413),
            .I(N__31391));
    InMux I__7173 (
            .O(N__31412),
            .I(N__31391));
    InMux I__7172 (
            .O(N__31411),
            .I(N__31386));
    InMux I__7171 (
            .O(N__31410),
            .I(N__31386));
    InMux I__7170 (
            .O(N__31409),
            .I(N__31381));
    InMux I__7169 (
            .O(N__31408),
            .I(N__31381));
    InMux I__7168 (
            .O(N__31407),
            .I(N__31378));
    InMux I__7167 (
            .O(N__31406),
            .I(N__31373));
    InMux I__7166 (
            .O(N__31405),
            .I(N__31373));
    InMux I__7165 (
            .O(N__31402),
            .I(N__31370));
    InMux I__7164 (
            .O(N__31401),
            .I(N__31365));
    InMux I__7163 (
            .O(N__31400),
            .I(N__31365));
    InMux I__7162 (
            .O(N__31399),
            .I(N__31362));
    Span4Mux_v I__7161 (
            .O(N__31396),
            .I(N__31355));
    LocalMux I__7160 (
            .O(N__31391),
            .I(N__31355));
    LocalMux I__7159 (
            .O(N__31386),
            .I(N__31355));
    LocalMux I__7158 (
            .O(N__31381),
            .I(N__31349));
    LocalMux I__7157 (
            .O(N__31378),
            .I(N__31346));
    LocalMux I__7156 (
            .O(N__31373),
            .I(N__31339));
    LocalMux I__7155 (
            .O(N__31370),
            .I(N__31339));
    LocalMux I__7154 (
            .O(N__31365),
            .I(N__31339));
    LocalMux I__7153 (
            .O(N__31362),
            .I(N__31336));
    Span4Mux_h I__7152 (
            .O(N__31355),
            .I(N__31333));
    CascadeMux I__7151 (
            .O(N__31354),
            .I(N__31330));
    InMux I__7150 (
            .O(N__31353),
            .I(N__31327));
    InMux I__7149 (
            .O(N__31352),
            .I(N__31324));
    Span4Mux_v I__7148 (
            .O(N__31349),
            .I(N__31321));
    Span4Mux_h I__7147 (
            .O(N__31346),
            .I(N__31316));
    Span4Mux_v I__7146 (
            .O(N__31339),
            .I(N__31316));
    Span4Mux_v I__7145 (
            .O(N__31336),
            .I(N__31311));
    Span4Mux_v I__7144 (
            .O(N__31333),
            .I(N__31311));
    InMux I__7143 (
            .O(N__31330),
            .I(N__31308));
    LocalMux I__7142 (
            .O(N__31327),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__7141 (
            .O(N__31324),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__7140 (
            .O(N__31321),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__7139 (
            .O(N__31316),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    Odrv4 I__7138 (
            .O(N__31311),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    LocalMux I__7137 (
            .O(N__31308),
            .I(\this_vga_signals.M_vcounter_qZ0Z_3 ));
    CascadeMux I__7136 (
            .O(N__31295),
            .I(N__31290));
    InMux I__7135 (
            .O(N__31294),
            .I(N__31281));
    InMux I__7134 (
            .O(N__31293),
            .I(N__31281));
    InMux I__7133 (
            .O(N__31290),
            .I(N__31278));
    InMux I__7132 (
            .O(N__31289),
            .I(N__31275));
    InMux I__7131 (
            .O(N__31288),
            .I(N__31269));
    InMux I__7130 (
            .O(N__31287),
            .I(N__31264));
    InMux I__7129 (
            .O(N__31286),
            .I(N__31264));
    LocalMux I__7128 (
            .O(N__31281),
            .I(N__31261));
    LocalMux I__7127 (
            .O(N__31278),
            .I(N__31257));
    LocalMux I__7126 (
            .O(N__31275),
            .I(N__31254));
    InMux I__7125 (
            .O(N__31274),
            .I(N__31249));
    InMux I__7124 (
            .O(N__31273),
            .I(N__31249));
    CascadeMux I__7123 (
            .O(N__31272),
            .I(N__31246));
    LocalMux I__7122 (
            .O(N__31269),
            .I(N__31243));
    LocalMux I__7121 (
            .O(N__31264),
            .I(N__31238));
    Span4Mux_h I__7120 (
            .O(N__31261),
            .I(N__31238));
    InMux I__7119 (
            .O(N__31260),
            .I(N__31235));
    Span4Mux_h I__7118 (
            .O(N__31257),
            .I(N__31230));
    Span4Mux_v I__7117 (
            .O(N__31254),
            .I(N__31230));
    LocalMux I__7116 (
            .O(N__31249),
            .I(N__31227));
    InMux I__7115 (
            .O(N__31246),
            .I(N__31223));
    Span4Mux_v I__7114 (
            .O(N__31243),
            .I(N__31220));
    Span4Mux_v I__7113 (
            .O(N__31238),
            .I(N__31217));
    LocalMux I__7112 (
            .O(N__31235),
            .I(N__31212));
    Span4Mux_v I__7111 (
            .O(N__31230),
            .I(N__31212));
    Span4Mux_v I__7110 (
            .O(N__31227),
            .I(N__31209));
    InMux I__7109 (
            .O(N__31226),
            .I(N__31206));
    LocalMux I__7108 (
            .O(N__31223),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__7107 (
            .O(N__31220),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__7106 (
            .O(N__31217),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__7105 (
            .O(N__31212),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    Odrv4 I__7104 (
            .O(N__31209),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    LocalMux I__7103 (
            .O(N__31206),
            .I(\this_vga_signals.M_vcounter_qZ0Z_2 ));
    InMux I__7102 (
            .O(N__31193),
            .I(N__31190));
    LocalMux I__7101 (
            .O(N__31190),
            .I(\this_vga_signals.N_5_i_1 ));
    InMux I__7100 (
            .O(N__31187),
            .I(N__31184));
    LocalMux I__7099 (
            .O(N__31184),
            .I(N__31181));
    Odrv12 I__7098 (
            .O(N__31181),
            .I(\this_vga_signals.N_5786_0_0 ));
    InMux I__7097 (
            .O(N__31178),
            .I(N__31175));
    LocalMux I__7096 (
            .O(N__31175),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ));
    CascadeMux I__7095 (
            .O(N__31172),
            .I(N__31169));
    InMux I__7094 (
            .O(N__31169),
            .I(N__31166));
    LocalMux I__7093 (
            .O(N__31166),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_x1 ));
    InMux I__7092 (
            .O(N__31163),
            .I(N__31160));
    LocalMux I__7091 (
            .O(N__31160),
            .I(N__31156));
    InMux I__7090 (
            .O(N__31159),
            .I(N__31153));
    Span4Mux_h I__7089 (
            .O(N__31156),
            .I(N__31150));
    LocalMux I__7088 (
            .O(N__31153),
            .I(\this_vga_signals.CO0_0_i_i ));
    Odrv4 I__7087 (
            .O(N__31150),
            .I(\this_vga_signals.CO0_0_i_i ));
    InMux I__7086 (
            .O(N__31145),
            .I(N__31142));
    LocalMux I__7085 (
            .O(N__31142),
            .I(N__31139));
    Span4Mux_h I__7084 (
            .O(N__31139),
            .I(N__31136));
    Odrv4 I__7083 (
            .O(N__31136),
            .I(\this_vga_signals.N_12_0 ));
    CascadeMux I__7082 (
            .O(N__31133),
            .I(\this_vga_signals.N_12_0_cascade_ ));
    InMux I__7081 (
            .O(N__31130),
            .I(N__31126));
    InMux I__7080 (
            .O(N__31129),
            .I(N__31123));
    LocalMux I__7079 (
            .O(N__31126),
            .I(N__31119));
    LocalMux I__7078 (
            .O(N__31123),
            .I(N__31116));
    InMux I__7077 (
            .O(N__31122),
            .I(N__31113));
    Span4Mux_v I__7076 (
            .O(N__31119),
            .I(N__31110));
    Odrv4 I__7075 (
            .O(N__31116),
            .I(\this_vga_signals.N_7_1_0 ));
    LocalMux I__7074 (
            .O(N__31113),
            .I(\this_vga_signals.N_7_1_0 ));
    Odrv4 I__7073 (
            .O(N__31110),
            .I(\this_vga_signals.N_7_1_0 ));
    InMux I__7072 (
            .O(N__31103),
            .I(N__31100));
    LocalMux I__7071 (
            .O(N__31100),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1 ));
    CascadeMux I__7070 (
            .O(N__31097),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_ ));
    InMux I__7069 (
            .O(N__31094),
            .I(N__31091));
    LocalMux I__7068 (
            .O(N__31091),
            .I(N__31088));
    Span4Mux_h I__7067 (
            .O(N__31088),
            .I(N__31085));
    Odrv4 I__7066 (
            .O(N__31085),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_0 ));
    InMux I__7065 (
            .O(N__31082),
            .I(N__31079));
    LocalMux I__7064 (
            .O(N__31079),
            .I(\this_vga_signals.g0_0_1 ));
    InMux I__7063 (
            .O(N__31076),
            .I(N__31073));
    LocalMux I__7062 (
            .O(N__31073),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_x0 ));
    CascadeMux I__7061 (
            .O(N__31070),
            .I(N__31066));
    CascadeMux I__7060 (
            .O(N__31069),
            .I(N__31061));
    InMux I__7059 (
            .O(N__31066),
            .I(N__31058));
    InMux I__7058 (
            .O(N__31065),
            .I(N__31053));
    InMux I__7057 (
            .O(N__31064),
            .I(N__31053));
    InMux I__7056 (
            .O(N__31061),
            .I(N__31050));
    LocalMux I__7055 (
            .O(N__31058),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_1 ));
    LocalMux I__7054 (
            .O(N__31053),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_1 ));
    LocalMux I__7053 (
            .O(N__31050),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_1 ));
    InMux I__7052 (
            .O(N__31043),
            .I(N__31040));
    LocalMux I__7051 (
            .O(N__31040),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ));
    InMux I__7050 (
            .O(N__31037),
            .I(N__31034));
    LocalMux I__7049 (
            .O(N__31034),
            .I(N__31030));
    InMux I__7048 (
            .O(N__31033),
            .I(N__31027));
    Span4Mux_h I__7047 (
            .O(N__31030),
            .I(N__31024));
    LocalMux I__7046 (
            .O(N__31027),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    Odrv4 I__7045 (
            .O(N__31024),
            .I(\this_vga_signals.mult1_un54_sum_axb1 ));
    CascadeMux I__7044 (
            .O(N__31019),
            .I(N__31008));
    CascadeMux I__7043 (
            .O(N__31018),
            .I(N__31005));
    CascadeMux I__7042 (
            .O(N__31017),
            .I(N__31002));
    CascadeMux I__7041 (
            .O(N__31016),
            .I(N__30999));
    CascadeMux I__7040 (
            .O(N__31015),
            .I(N__30996));
    InMux I__7039 (
            .O(N__31014),
            .I(N__30992));
    IoInMux I__7038 (
            .O(N__31013),
            .I(N__30980));
    InMux I__7037 (
            .O(N__31012),
            .I(N__30977));
    InMux I__7036 (
            .O(N__31011),
            .I(N__30972));
    InMux I__7035 (
            .O(N__31008),
            .I(N__30972));
    InMux I__7034 (
            .O(N__31005),
            .I(N__30967));
    InMux I__7033 (
            .O(N__31002),
            .I(N__30967));
    InMux I__7032 (
            .O(N__30999),
            .I(N__30960));
    InMux I__7031 (
            .O(N__30996),
            .I(N__30960));
    InMux I__7030 (
            .O(N__30995),
            .I(N__30960));
    LocalMux I__7029 (
            .O(N__30992),
            .I(N__30957));
    InMux I__7028 (
            .O(N__30991),
            .I(N__30954));
    InMux I__7027 (
            .O(N__30990),
            .I(N__30951));
    InMux I__7026 (
            .O(N__30989),
            .I(N__30946));
    InMux I__7025 (
            .O(N__30988),
            .I(N__30946));
    InMux I__7024 (
            .O(N__30987),
            .I(N__30939));
    InMux I__7023 (
            .O(N__30986),
            .I(N__30939));
    InMux I__7022 (
            .O(N__30985),
            .I(N__30939));
    InMux I__7021 (
            .O(N__30984),
            .I(N__30936));
    InMux I__7020 (
            .O(N__30983),
            .I(N__30933));
    LocalMux I__7019 (
            .O(N__30980),
            .I(N__30929));
    LocalMux I__7018 (
            .O(N__30977),
            .I(N__30926));
    LocalMux I__7017 (
            .O(N__30972),
            .I(N__30915));
    LocalMux I__7016 (
            .O(N__30967),
            .I(N__30915));
    LocalMux I__7015 (
            .O(N__30960),
            .I(N__30915));
    Span4Mux_h I__7014 (
            .O(N__30957),
            .I(N__30915));
    LocalMux I__7013 (
            .O(N__30954),
            .I(N__30915));
    LocalMux I__7012 (
            .O(N__30951),
            .I(N__30912));
    LocalMux I__7011 (
            .O(N__30946),
            .I(N__30909));
    LocalMux I__7010 (
            .O(N__30939),
            .I(N__30906));
    LocalMux I__7009 (
            .O(N__30936),
            .I(N__30901));
    LocalMux I__7008 (
            .O(N__30933),
            .I(N__30901));
    CascadeMux I__7007 (
            .O(N__30932),
            .I(N__30896));
    IoSpan4Mux I__7006 (
            .O(N__30929),
            .I(N__30891));
    Span4Mux_h I__7005 (
            .O(N__30926),
            .I(N__30884));
    Span4Mux_h I__7004 (
            .O(N__30915),
            .I(N__30884));
    Span4Mux_v I__7003 (
            .O(N__30912),
            .I(N__30884));
    Span4Mux_v I__7002 (
            .O(N__30909),
            .I(N__30881));
    Span4Mux_v I__7001 (
            .O(N__30906),
            .I(N__30878));
    Span4Mux_h I__7000 (
            .O(N__30901),
            .I(N__30875));
    InMux I__6999 (
            .O(N__30900),
            .I(N__30870));
    InMux I__6998 (
            .O(N__30899),
            .I(N__30870));
    InMux I__6997 (
            .O(N__30896),
            .I(N__30863));
    InMux I__6996 (
            .O(N__30895),
            .I(N__30863));
    InMux I__6995 (
            .O(N__30894),
            .I(N__30863));
    IoSpan4Mux I__6994 (
            .O(N__30891),
            .I(N__30860));
    Span4Mux_v I__6993 (
            .O(N__30884),
            .I(N__30857));
    Span4Mux_h I__6992 (
            .O(N__30881),
            .I(N__30852));
    Span4Mux_h I__6991 (
            .O(N__30878),
            .I(N__30852));
    Span4Mux_v I__6990 (
            .O(N__30875),
            .I(N__30849));
    LocalMux I__6989 (
            .O(N__30870),
            .I(N__30844));
    LocalMux I__6988 (
            .O(N__30863),
            .I(N__30844));
    Sp12to4 I__6987 (
            .O(N__30860),
            .I(N__30841));
    Span4Mux_h I__6986 (
            .O(N__30857),
            .I(N__30838));
    Span4Mux_h I__6985 (
            .O(N__30852),
            .I(N__30835));
    Span4Mux_v I__6984 (
            .O(N__30849),
            .I(N__30832));
    Span12Mux_v I__6983 (
            .O(N__30844),
            .I(N__30827));
    Span12Mux_s9_h I__6982 (
            .O(N__30841),
            .I(N__30827));
    Odrv4 I__6981 (
            .O(N__30838),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__6980 (
            .O(N__30835),
            .I(M_this_reset_cond_out_0));
    Odrv4 I__6979 (
            .O(N__30832),
            .I(M_this_reset_cond_out_0));
    Odrv12 I__6978 (
            .O(N__30827),
            .I(M_this_reset_cond_out_0));
    InMux I__6977 (
            .O(N__30818),
            .I(N__30809));
    InMux I__6976 (
            .O(N__30817),
            .I(N__30809));
    InMux I__6975 (
            .O(N__30816),
            .I(N__30802));
    InMux I__6974 (
            .O(N__30815),
            .I(N__30802));
    InMux I__6973 (
            .O(N__30814),
            .I(N__30802));
    LocalMux I__6972 (
            .O(N__30809),
            .I(N__30795));
    LocalMux I__6971 (
            .O(N__30802),
            .I(N__30792));
    InMux I__6970 (
            .O(N__30801),
            .I(N__30789));
    InMux I__6969 (
            .O(N__30800),
            .I(N__30782));
    InMux I__6968 (
            .O(N__30799),
            .I(N__30782));
    InMux I__6967 (
            .O(N__30798),
            .I(N__30782));
    Span4Mux_v I__6966 (
            .O(N__30795),
            .I(N__30778));
    Span4Mux_v I__6965 (
            .O(N__30792),
            .I(N__30775));
    LocalMux I__6964 (
            .O(N__30789),
            .I(N__30772));
    LocalMux I__6963 (
            .O(N__30782),
            .I(N__30769));
    InMux I__6962 (
            .O(N__30781),
            .I(N__30766));
    Sp12to4 I__6961 (
            .O(N__30778),
            .I(N__30763));
    Sp12to4 I__6960 (
            .O(N__30775),
            .I(N__30760));
    Span4Mux_h I__6959 (
            .O(N__30772),
            .I(N__30757));
    Span4Mux_h I__6958 (
            .O(N__30769),
            .I(N__30752));
    LocalMux I__6957 (
            .O(N__30766),
            .I(N__30752));
    Span12Mux_h I__6956 (
            .O(N__30763),
            .I(N__30743));
    Span12Mux_h I__6955 (
            .O(N__30760),
            .I(N__30743));
    Sp12to4 I__6954 (
            .O(N__30757),
            .I(N__30743));
    Sp12to4 I__6953 (
            .O(N__30752),
            .I(N__30743));
    Span12Mux_v I__6952 (
            .O(N__30743),
            .I(N__30740));
    Span12Mux_v I__6951 (
            .O(N__30740),
            .I(N__30737));
    Odrv12 I__6950 (
            .O(N__30737),
            .I(rst_n_c));
    InMux I__6949 (
            .O(N__30734),
            .I(N__30731));
    LocalMux I__6948 (
            .O(N__30731),
            .I(\this_reset_cond.M_stage_qZ0Z_7 ));
    InMux I__6947 (
            .O(N__30728),
            .I(N__30725));
    LocalMux I__6946 (
            .O(N__30725),
            .I(\this_reset_cond.M_stage_qZ0Z_8 ));
    CEMux I__6945 (
            .O(N__30722),
            .I(N__30719));
    LocalMux I__6944 (
            .O(N__30719),
            .I(N__30715));
    CEMux I__6943 (
            .O(N__30718),
            .I(N__30712));
    Span4Mux_h I__6942 (
            .O(N__30715),
            .I(N__30709));
    LocalMux I__6941 (
            .O(N__30712),
            .I(N__30706));
    Span4Mux_v I__6940 (
            .O(N__30709),
            .I(N__30703));
    Span4Mux_h I__6939 (
            .O(N__30706),
            .I(N__30700));
    Span4Mux_h I__6938 (
            .O(N__30703),
            .I(N__30697));
    Span4Mux_h I__6937 (
            .O(N__30700),
            .I(N__30694));
    Odrv4 I__6936 (
            .O(N__30697),
            .I(\this_spr_ram.mem_WE_10 ));
    Odrv4 I__6935 (
            .O(N__30694),
            .I(\this_spr_ram.mem_WE_10 ));
    InMux I__6934 (
            .O(N__30689),
            .I(N__30686));
    LocalMux I__6933 (
            .O(N__30686),
            .I(\this_vga_signals.N_12_0_0 ));
    CascadeMux I__6932 (
            .O(N__30683),
            .I(N__30680));
    InMux I__6931 (
            .O(N__30680),
            .I(N__30677));
    LocalMux I__6930 (
            .O(N__30677),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ));
    InMux I__6929 (
            .O(N__30674),
            .I(N__30671));
    LocalMux I__6928 (
            .O(N__30671),
            .I(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ));
    CascadeMux I__6927 (
            .O(N__30668),
            .I(\this_vga_signals.vaddress_c2_cascade_ ));
    InMux I__6926 (
            .O(N__30665),
            .I(N__30662));
    LocalMux I__6925 (
            .O(N__30662),
            .I(N__30659));
    Odrv4 I__6924 (
            .O(N__30659),
            .I(\this_vga_signals.g1_1 ));
    InMux I__6923 (
            .O(N__30656),
            .I(N__30653));
    LocalMux I__6922 (
            .O(N__30653),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_0 ));
    CascadeMux I__6921 (
            .O(N__30650),
            .I(\this_vga_signals.g0_1_0_cascade_ ));
    InMux I__6920 (
            .O(N__30647),
            .I(N__30644));
    LocalMux I__6919 (
            .O(N__30644),
            .I(N__30641));
    Odrv12 I__6918 (
            .O(N__30641),
            .I(\this_vga_signals.N_7_1_0_2 ));
    CascadeMux I__6917 (
            .O(N__30638),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ));
    CascadeMux I__6916 (
            .O(N__30635),
            .I(N__30632));
    InMux I__6915 (
            .O(N__30632),
            .I(N__30629));
    LocalMux I__6914 (
            .O(N__30629),
            .I(N__30626));
    Odrv4 I__6913 (
            .O(N__30626),
            .I(\this_vga_signals.g3_1 ));
    InMux I__6912 (
            .O(N__30623),
            .I(N__30620));
    LocalMux I__6911 (
            .O(N__30620),
            .I(N__30616));
    InMux I__6910 (
            .O(N__30619),
            .I(N__30613));
    Span4Mux_h I__6909 (
            .O(N__30616),
            .I(N__30610));
    LocalMux I__6908 (
            .O(N__30613),
            .I(N__30607));
    Odrv4 I__6907 (
            .O(N__30610),
            .I(\this_vga_signals.g1_3 ));
    Odrv12 I__6906 (
            .O(N__30607),
            .I(\this_vga_signals.g1_3 ));
    InMux I__6905 (
            .O(N__30602),
            .I(N__30599));
    LocalMux I__6904 (
            .O(N__30599),
            .I(\this_vga_signals.N_7_1_0_0 ));
    InMux I__6903 (
            .O(N__30596),
            .I(N__30593));
    LocalMux I__6902 (
            .O(N__30593),
            .I(\this_vga_signals.g0_1_0_0 ));
    InMux I__6901 (
            .O(N__30590),
            .I(N__30587));
    LocalMux I__6900 (
            .O(N__30587),
            .I(N__30584));
    Span4Mux_v I__6899 (
            .O(N__30584),
            .I(N__30577));
    InMux I__6898 (
            .O(N__30583),
            .I(N__30572));
    InMux I__6897 (
            .O(N__30582),
            .I(N__30572));
    InMux I__6896 (
            .O(N__30581),
            .I(N__30569));
    InMux I__6895 (
            .O(N__30580),
            .I(N__30566));
    Span4Mux_h I__6894 (
            .O(N__30577),
            .I(N__30554));
    LocalMux I__6893 (
            .O(N__30572),
            .I(N__30551));
    LocalMux I__6892 (
            .O(N__30569),
            .I(N__30548));
    LocalMux I__6891 (
            .O(N__30566),
            .I(N__30545));
    InMux I__6890 (
            .O(N__30565),
            .I(N__30538));
    InMux I__6889 (
            .O(N__30564),
            .I(N__30538));
    InMux I__6888 (
            .O(N__30563),
            .I(N__30538));
    InMux I__6887 (
            .O(N__30562),
            .I(N__30531));
    InMux I__6886 (
            .O(N__30561),
            .I(N__30531));
    InMux I__6885 (
            .O(N__30560),
            .I(N__30531));
    InMux I__6884 (
            .O(N__30559),
            .I(N__30524));
    InMux I__6883 (
            .O(N__30558),
            .I(N__30524));
    InMux I__6882 (
            .O(N__30557),
            .I(N__30524));
    Odrv4 I__6881 (
            .O(N__30554),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    Odrv4 I__6880 (
            .O(N__30551),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    Odrv4 I__6879 (
            .O(N__30548),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    Odrv4 I__6878 (
            .O(N__30545),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__6877 (
            .O(N__30538),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__6876 (
            .O(N__30531),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    LocalMux I__6875 (
            .O(N__30524),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns ));
    InMux I__6874 (
            .O(N__30509),
            .I(N__30506));
    LocalMux I__6873 (
            .O(N__30506),
            .I(\this_vga_signals.g1_0 ));
    CascadeMux I__6872 (
            .O(N__30503),
            .I(N__30495));
    CascadeMux I__6871 (
            .O(N__30502),
            .I(N__30492));
    InMux I__6870 (
            .O(N__30501),
            .I(N__30489));
    InMux I__6869 (
            .O(N__30500),
            .I(N__30481));
    InMux I__6868 (
            .O(N__30499),
            .I(N__30481));
    CascadeMux I__6867 (
            .O(N__30498),
            .I(N__30478));
    InMux I__6866 (
            .O(N__30495),
            .I(N__30475));
    InMux I__6865 (
            .O(N__30492),
            .I(N__30472));
    LocalMux I__6864 (
            .O(N__30489),
            .I(N__30469));
    InMux I__6863 (
            .O(N__30488),
            .I(N__30466));
    CascadeMux I__6862 (
            .O(N__30487),
            .I(N__30463));
    CascadeMux I__6861 (
            .O(N__30486),
            .I(N__30460));
    LocalMux I__6860 (
            .O(N__30481),
            .I(N__30457));
    InMux I__6859 (
            .O(N__30478),
            .I(N__30454));
    LocalMux I__6858 (
            .O(N__30475),
            .I(N__30449));
    LocalMux I__6857 (
            .O(N__30472),
            .I(N__30449));
    Span4Mux_v I__6856 (
            .O(N__30469),
            .I(N__30444));
    LocalMux I__6855 (
            .O(N__30466),
            .I(N__30444));
    InMux I__6854 (
            .O(N__30463),
            .I(N__30439));
    InMux I__6853 (
            .O(N__30460),
            .I(N__30439));
    Odrv12 I__6852 (
            .O(N__30457),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6851 (
            .O(N__30454),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    Odrv4 I__6850 (
            .O(N__30449),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    Odrv4 I__6849 (
            .O(N__30444),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    LocalMux I__6848 (
            .O(N__30439),
            .I(\this_vga_signals.mult1_un54_sum_c2_0 ));
    InMux I__6847 (
            .O(N__30428),
            .I(N__30425));
    LocalMux I__6846 (
            .O(N__30425),
            .I(\this_vga_signals.g0_29_1 ));
    CascadeMux I__6845 (
            .O(N__30422),
            .I(\this_vga_signals.g1_0_cascade_ ));
    CascadeMux I__6844 (
            .O(N__30419),
            .I(N__30414));
    InMux I__6843 (
            .O(N__30418),
            .I(N__30409));
    InMux I__6842 (
            .O(N__30417),
            .I(N__30404));
    InMux I__6841 (
            .O(N__30414),
            .I(N__30404));
    CascadeMux I__6840 (
            .O(N__30413),
            .I(N__30400));
    CascadeMux I__6839 (
            .O(N__30412),
            .I(N__30394));
    LocalMux I__6838 (
            .O(N__30409),
            .I(N__30389));
    LocalMux I__6837 (
            .O(N__30404),
            .I(N__30386));
    InMux I__6836 (
            .O(N__30403),
            .I(N__30383));
    InMux I__6835 (
            .O(N__30400),
            .I(N__30378));
    InMux I__6834 (
            .O(N__30399),
            .I(N__30378));
    InMux I__6833 (
            .O(N__30398),
            .I(N__30371));
    InMux I__6832 (
            .O(N__30397),
            .I(N__30371));
    InMux I__6831 (
            .O(N__30394),
            .I(N__30371));
    InMux I__6830 (
            .O(N__30393),
            .I(N__30366));
    InMux I__6829 (
            .O(N__30392),
            .I(N__30366));
    Odrv4 I__6828 (
            .O(N__30389),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    Odrv4 I__6827 (
            .O(N__30386),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    LocalMux I__6826 (
            .O(N__30383),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    LocalMux I__6825 (
            .O(N__30378),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    LocalMux I__6824 (
            .O(N__30371),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    LocalMux I__6823 (
            .O(N__30366),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0));
    InMux I__6822 (
            .O(N__30353),
            .I(N__30350));
    LocalMux I__6821 (
            .O(N__30350),
            .I(\this_vga_signals.g0_3 ));
    InMux I__6820 (
            .O(N__30347),
            .I(N__30344));
    LocalMux I__6819 (
            .O(N__30344),
            .I(N__30341));
    Odrv4 I__6818 (
            .O(N__30341),
            .I(\this_reset_cond.M_stage_qZ0Z_6 ));
    CascadeMux I__6817 (
            .O(N__30338),
            .I(N__30335));
    InMux I__6816 (
            .O(N__30335),
            .I(N__30332));
    LocalMux I__6815 (
            .O(N__30332),
            .I(N__30329));
    Odrv4 I__6814 (
            .O(N__30329),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4 ));
    CascadeMux I__6813 (
            .O(N__30326),
            .I(\this_vga_signals.g0_2_0_0_cascade_ ));
    InMux I__6812 (
            .O(N__30323),
            .I(N__30320));
    LocalMux I__6811 (
            .O(N__30320),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_4 ));
    InMux I__6810 (
            .O(N__30317),
            .I(N__30314));
    LocalMux I__6809 (
            .O(N__30314),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0 ));
    CascadeMux I__6808 (
            .O(N__30311),
            .I(N__30308));
    InMux I__6807 (
            .O(N__30308),
            .I(N__30305));
    LocalMux I__6806 (
            .O(N__30305),
            .I(\this_vga_signals.g0_6_0 ));
    CascadeMux I__6805 (
            .O(N__30302),
            .I(N__30299));
    InMux I__6804 (
            .O(N__30299),
            .I(N__30296));
    LocalMux I__6803 (
            .O(N__30296),
            .I(\this_vga_signals.g0_0_0_1 ));
    InMux I__6802 (
            .O(N__30293),
            .I(N__30290));
    LocalMux I__6801 (
            .O(N__30290),
            .I(\this_vga_signals.g0_5_5_N_2L1 ));
    CascadeMux I__6800 (
            .O(N__30287),
            .I(N__30284));
    InMux I__6799 (
            .O(N__30284),
            .I(N__30272));
    InMux I__6798 (
            .O(N__30283),
            .I(N__30269));
    InMux I__6797 (
            .O(N__30282),
            .I(N__30266));
    InMux I__6796 (
            .O(N__30281),
            .I(N__30261));
    InMux I__6795 (
            .O(N__30280),
            .I(N__30261));
    InMux I__6794 (
            .O(N__30279),
            .I(N__30254));
    InMux I__6793 (
            .O(N__30278),
            .I(N__30254));
    InMux I__6792 (
            .O(N__30277),
            .I(N__30254));
    InMux I__6791 (
            .O(N__30276),
            .I(N__30249));
    InMux I__6790 (
            .O(N__30275),
            .I(N__30249));
    LocalMux I__6789 (
            .O(N__30272),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    LocalMux I__6788 (
            .O(N__30269),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    LocalMux I__6787 (
            .O(N__30266),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    LocalMux I__6786 (
            .O(N__30261),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    LocalMux I__6785 (
            .O(N__30254),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    LocalMux I__6784 (
            .O(N__30249),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0));
    InMux I__6783 (
            .O(N__30236),
            .I(N__30233));
    LocalMux I__6782 (
            .O(N__30233),
            .I(\this_vga_signals.g0_5_0 ));
    CascadeMux I__6781 (
            .O(N__30230),
            .I(N__30224));
    InMux I__6780 (
            .O(N__30229),
            .I(N__30214));
    InMux I__6779 (
            .O(N__30228),
            .I(N__30214));
    InMux I__6778 (
            .O(N__30227),
            .I(N__30211));
    InMux I__6777 (
            .O(N__30224),
            .I(N__30204));
    InMux I__6776 (
            .O(N__30223),
            .I(N__30204));
    InMux I__6775 (
            .O(N__30222),
            .I(N__30204));
    InMux I__6774 (
            .O(N__30221),
            .I(N__30197));
    InMux I__6773 (
            .O(N__30220),
            .I(N__30197));
    InMux I__6772 (
            .O(N__30219),
            .I(N__30197));
    LocalMux I__6771 (
            .O(N__30214),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__6770 (
            .O(N__30211),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__6769 (
            .O(N__30204),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    LocalMux I__6768 (
            .O(N__30197),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3 ));
    CascadeMux I__6767 (
            .O(N__30188),
            .I(\this_vga_signals.mult1_un54_sum_c2_0_cascade_ ));
    CascadeMux I__6766 (
            .O(N__30185),
            .I(\this_vga_signals.g1_1_0_0_cascade_ ));
    InMux I__6765 (
            .O(N__30182),
            .I(N__30179));
    LocalMux I__6764 (
            .O(N__30179),
            .I(\this_vga_signals.N_20_0 ));
    CascadeMux I__6763 (
            .O(N__30176),
            .I(\this_vga_signals.g0_2_0_3_cascade_ ));
    InMux I__6762 (
            .O(N__30173),
            .I(N__30170));
    LocalMux I__6761 (
            .O(N__30170),
            .I(\this_vga_signals.g0_0_0_1_0 ));
    InMux I__6760 (
            .O(N__30167),
            .I(N__30164));
    LocalMux I__6759 (
            .O(N__30164),
            .I(\this_vga_signals.g0_0_0 ));
    CascadeMux I__6758 (
            .O(N__30161),
            .I(\this_vga_signals.vaddress_c5_a0_0_cascade_ ));
    CascadeMux I__6757 (
            .O(N__30158),
            .I(\this_vga_signals.vaddress_9_cascade_ ));
    CascadeMux I__6756 (
            .O(N__30155),
            .I(\this_vga_signals.g1_3_0_cascade_ ));
    CascadeMux I__6755 (
            .O(N__30152),
            .I(\this_vga_signals.N_5_0_cascade_ ));
    CascadeMux I__6754 (
            .O(N__30149),
            .I(N__30146));
    InMux I__6753 (
            .O(N__30146),
            .I(N__30143));
    LocalMux I__6752 (
            .O(N__30143),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_0_0 ));
    InMux I__6751 (
            .O(N__30140),
            .I(N__30137));
    LocalMux I__6750 (
            .O(N__30137),
            .I(\this_vga_signals.N_4_1 ));
    CascadeMux I__6749 (
            .O(N__30134),
            .I(\this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_ ));
    InMux I__6748 (
            .O(N__30131),
            .I(N__30128));
    LocalMux I__6747 (
            .O(N__30128),
            .I(\this_vga_signals.mult1_un54_sum_c3_x1 ));
    IoInMux I__6746 (
            .O(N__30125),
            .I(N__30122));
    LocalMux I__6745 (
            .O(N__30122),
            .I(N__30119));
    Span4Mux_s2_v I__6744 (
            .O(N__30119),
            .I(N__30116));
    Odrv4 I__6743 (
            .O(N__30116),
            .I(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO));
    CEMux I__6742 (
            .O(N__30113),
            .I(N__30110));
    LocalMux I__6741 (
            .O(N__30110),
            .I(N__30106));
    CEMux I__6740 (
            .O(N__30109),
            .I(N__30103));
    Span4Mux_v I__6739 (
            .O(N__30106),
            .I(N__30100));
    LocalMux I__6738 (
            .O(N__30103),
            .I(N__30097));
    Span4Mux_h I__6737 (
            .O(N__30100),
            .I(N__30092));
    Span4Mux_h I__6736 (
            .O(N__30097),
            .I(N__30092));
    Span4Mux_h I__6735 (
            .O(N__30092),
            .I(N__30089));
    Odrv4 I__6734 (
            .O(N__30089),
            .I(\this_spr_ram.mem_WE_8 ));
    InMux I__6733 (
            .O(N__30086),
            .I(N__30083));
    LocalMux I__6732 (
            .O(N__30083),
            .I(\this_vga_signals.m43_4 ));
    CascadeMux I__6731 (
            .O(N__30080),
            .I(N__30077));
    InMux I__6730 (
            .O(N__30077),
            .I(N__30074));
    LocalMux I__6729 (
            .O(N__30074),
            .I(\this_vga_signals.vaddress_c3_d_0 ));
    InMux I__6728 (
            .O(N__30071),
            .I(N__30068));
    LocalMux I__6727 (
            .O(N__30068),
            .I(N__30065));
    Span4Mux_v I__6726 (
            .O(N__30065),
            .I(N__30062));
    Odrv4 I__6725 (
            .O(N__30062),
            .I(\this_vga_signals.g0_1_0_1 ));
    CascadeMux I__6724 (
            .O(N__30059),
            .I(\this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_ ));
    CascadeMux I__6723 (
            .O(N__30056),
            .I(\this_vga_signals.CO0_0_i_i_cascade_ ));
    CascadeMux I__6722 (
            .O(N__30053),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_ ));
    CascadeMux I__6721 (
            .O(N__30050),
            .I(\this_vga_signals.N_5_i_0_cascade_ ));
    InMux I__6720 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__6719 (
            .O(N__30044),
            .I(N__30041));
    Odrv4 I__6718 (
            .O(N__30041),
            .I(\this_vga_signals.g1_0_0 ));
    CascadeMux I__6717 (
            .O(N__30038),
            .I(N__30035));
    InMux I__6716 (
            .O(N__30035),
            .I(N__30032));
    LocalMux I__6715 (
            .O(N__30032),
            .I(N__30029));
    Odrv4 I__6714 (
            .O(N__30029),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9 ));
    InMux I__6713 (
            .O(N__30026),
            .I(N__30023));
    LocalMux I__6712 (
            .O(N__30023),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2 ));
    CascadeMux I__6711 (
            .O(N__30020),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ));
    CascadeMux I__6710 (
            .O(N__30017),
            .I(N__30014));
    InMux I__6709 (
            .O(N__30014),
            .I(N__30011));
    LocalMux I__6708 (
            .O(N__30011),
            .I(\this_vga_signals.g0_i_x2_1 ));
    CascadeMux I__6707 (
            .O(N__30008),
            .I(\this_vga_signals.mult1_un54_sum_c3_x0_cascade_ ));
    CascadeMux I__6706 (
            .O(N__30005),
            .I(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_));
    InMux I__6705 (
            .O(N__30002),
            .I(N__29999));
    LocalMux I__6704 (
            .O(N__29999),
            .I(\this_vga_signals.g0_41_N_4L5_1 ));
    InMux I__6703 (
            .O(N__29996),
            .I(N__29993));
    LocalMux I__6702 (
            .O(N__29993),
            .I(N_6_i));
    CascadeMux I__6701 (
            .O(N__29990),
            .I(\this_vga_signals.g0_1_1_cascade_ ));
    InMux I__6700 (
            .O(N__29987),
            .I(N__29984));
    LocalMux I__6699 (
            .O(N__29984),
            .I(\this_vga_signals.mult1_un61_sum_c2_0_0 ));
    InMux I__6698 (
            .O(N__29981),
            .I(N__29978));
    LocalMux I__6697 (
            .O(N__29978),
            .I(\this_vga_signals.g1_4 ));
    InMux I__6696 (
            .O(N__29975),
            .I(N__29972));
    LocalMux I__6695 (
            .O(N__29972),
            .I(\this_vga_signals.g1_0_0_0 ));
    CascadeMux I__6694 (
            .O(N__29969),
            .I(\this_vga_signals.g1_0_1_0_cascade_ ));
    InMux I__6693 (
            .O(N__29966),
            .I(N__29963));
    LocalMux I__6692 (
            .O(N__29963),
            .I(\this_vga_signals.N_10 ));
    InMux I__6691 (
            .O(N__29960),
            .I(N__29957));
    LocalMux I__6690 (
            .O(N__29957),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_d_2_0 ));
    InMux I__6689 (
            .O(N__29954),
            .I(N__29951));
    LocalMux I__6688 (
            .O(N__29951),
            .I(\this_vga_signals.g0_0_i_0_1 ));
    CascadeMux I__6687 (
            .O(N__29948),
            .I(\this_vga_signals.N_10_i_cascade_ ));
    InMux I__6686 (
            .O(N__29945),
            .I(N__29942));
    LocalMux I__6685 (
            .O(N__29942),
            .I(N__29939));
    Span4Mux_h I__6684 (
            .O(N__29939),
            .I(N__29936));
    Odrv4 I__6683 (
            .O(N__29936),
            .I(\this_vga_signals.g2_1_2 ));
    InMux I__6682 (
            .O(N__29933),
            .I(N__29930));
    LocalMux I__6681 (
            .O(N__29930),
            .I(\this_vga_signals.N_10_i_0 ));
    CascadeMux I__6680 (
            .O(N__29927),
            .I(\this_vga_signals.g0_0_i_0_cascade_ ));
    InMux I__6679 (
            .O(N__29924),
            .I(N__29921));
    LocalMux I__6678 (
            .O(N__29921),
            .I(\this_vga_signals.if_m5_i_0_0 ));
    InMux I__6677 (
            .O(N__29918),
            .I(N__29915));
    LocalMux I__6676 (
            .O(N__29915),
            .I(\this_vga_signals.mult1_un68_sum_c3_0_0_0 ));
    InMux I__6675 (
            .O(N__29912),
            .I(N__29909));
    LocalMux I__6674 (
            .O(N__29909),
            .I(\this_vga_signals.if_N_10_0_0_0 ));
    InMux I__6673 (
            .O(N__29906),
            .I(N__29903));
    LocalMux I__6672 (
            .O(N__29903),
            .I(\this_vga_signals.g0_1_0_3 ));
    InMux I__6671 (
            .O(N__29900),
            .I(N__29897));
    LocalMux I__6670 (
            .O(N__29897),
            .I(\this_vga_signals.g0_1_1_0 ));
    CascadeMux I__6669 (
            .O(N__29894),
            .I(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ));
    InMux I__6668 (
            .O(N__29891),
            .I(N__29888));
    LocalMux I__6667 (
            .O(N__29888),
            .I(\this_vga_signals.g0_41_N_3L3_1 ));
    InMux I__6666 (
            .O(N__29885),
            .I(N__29882));
    LocalMux I__6665 (
            .O(N__29882),
            .I(\this_vga_signals.m43_5 ));
    IoInMux I__6664 (
            .O(N__29879),
            .I(N__29876));
    LocalMux I__6663 (
            .O(N__29876),
            .I(N__29873));
    Span4Mux_s3_v I__6662 (
            .O(N__29873),
            .I(N__29870));
    Span4Mux_h I__6661 (
            .O(N__29870),
            .I(N__29867));
    Span4Mux_v I__6660 (
            .O(N__29867),
            .I(N__29864));
    Sp12to4 I__6659 (
            .O(N__29864),
            .I(N__29861));
    Span12Mux_h I__6658 (
            .O(N__29861),
            .I(N__29858));
    Odrv12 I__6657 (
            .O(N__29858),
            .I(this_vga_signals_vsync_1_i));
    InMux I__6656 (
            .O(N__29855),
            .I(N__29852));
    LocalMux I__6655 (
            .O(N__29852),
            .I(N__29849));
    Span4Mux_v I__6654 (
            .O(N__29849),
            .I(N__29844));
    InMux I__6653 (
            .O(N__29848),
            .I(N__29841));
    InMux I__6652 (
            .O(N__29847),
            .I(N__29838));
    Span4Mux_h I__6651 (
            .O(N__29844),
            .I(N__29833));
    LocalMux I__6650 (
            .O(N__29841),
            .I(N__29833));
    LocalMux I__6649 (
            .O(N__29838),
            .I(N_52_0));
    Odrv4 I__6648 (
            .O(N__29833),
            .I(N_52_0));
    InMux I__6647 (
            .O(N__29828),
            .I(N__29825));
    LocalMux I__6646 (
            .O(N__29825),
            .I(N__29822));
    Span4Mux_h I__6645 (
            .O(N__29822),
            .I(N__29818));
    InMux I__6644 (
            .O(N__29821),
            .I(N__29815));
    Odrv4 I__6643 (
            .O(N__29818),
            .I(N_58_0));
    LocalMux I__6642 (
            .O(N__29815),
            .I(N_58_0));
    InMux I__6641 (
            .O(N__29810),
            .I(N__29806));
    InMux I__6640 (
            .O(N__29809),
            .I(N__29803));
    LocalMux I__6639 (
            .O(N__29806),
            .I(N__29798));
    LocalMux I__6638 (
            .O(N__29803),
            .I(N__29798));
    Span4Mux_v I__6637 (
            .O(N__29798),
            .I(N__29795));
    Odrv4 I__6636 (
            .O(N__29795),
            .I(\this_ppu.line_clk.M_last_qZ0 ));
    CEMux I__6635 (
            .O(N__29792),
            .I(N__29780));
    CascadeMux I__6634 (
            .O(N__29791),
            .I(N__29775));
    InMux I__6633 (
            .O(N__29790),
            .I(N__29767));
    InMux I__6632 (
            .O(N__29789),
            .I(N__29759));
    InMux I__6631 (
            .O(N__29788),
            .I(N__29759));
    InMux I__6630 (
            .O(N__29787),
            .I(N__29759));
    InMux I__6629 (
            .O(N__29786),
            .I(N__29750));
    InMux I__6628 (
            .O(N__29785),
            .I(N__29750));
    InMux I__6627 (
            .O(N__29784),
            .I(N__29750));
    InMux I__6626 (
            .O(N__29783),
            .I(N__29750));
    LocalMux I__6625 (
            .O(N__29780),
            .I(N__29747));
    CascadeMux I__6624 (
            .O(N__29779),
            .I(N__29744));
    InMux I__6623 (
            .O(N__29778),
            .I(N__29738));
    InMux I__6622 (
            .O(N__29775),
            .I(N__29738));
    InMux I__6621 (
            .O(N__29774),
            .I(N__29735));
    InMux I__6620 (
            .O(N__29773),
            .I(N__29726));
    InMux I__6619 (
            .O(N__29772),
            .I(N__29726));
    InMux I__6618 (
            .O(N__29771),
            .I(N__29721));
    InMux I__6617 (
            .O(N__29770),
            .I(N__29721));
    LocalMux I__6616 (
            .O(N__29767),
            .I(N__29718));
    InMux I__6615 (
            .O(N__29766),
            .I(N__29715));
    LocalMux I__6614 (
            .O(N__29759),
            .I(N__29712));
    LocalMux I__6613 (
            .O(N__29750),
            .I(N__29707));
    Span4Mux_h I__6612 (
            .O(N__29747),
            .I(N__29707));
    InMux I__6611 (
            .O(N__29744),
            .I(N__29702));
    InMux I__6610 (
            .O(N__29743),
            .I(N__29702));
    LocalMux I__6609 (
            .O(N__29738),
            .I(N__29699));
    LocalMux I__6608 (
            .O(N__29735),
            .I(N__29696));
    InMux I__6607 (
            .O(N__29734),
            .I(N__29687));
    InMux I__6606 (
            .O(N__29733),
            .I(N__29687));
    InMux I__6605 (
            .O(N__29732),
            .I(N__29687));
    InMux I__6604 (
            .O(N__29731),
            .I(N__29687));
    LocalMux I__6603 (
            .O(N__29726),
            .I(N__29678));
    LocalMux I__6602 (
            .O(N__29721),
            .I(N__29678));
    Span4Mux_v I__6601 (
            .O(N__29718),
            .I(N__29678));
    LocalMux I__6600 (
            .O(N__29715),
            .I(N__29678));
    Span4Mux_v I__6599 (
            .O(N__29712),
            .I(N__29673));
    Span4Mux_v I__6598 (
            .O(N__29707),
            .I(N__29673));
    LocalMux I__6597 (
            .O(N__29702),
            .I(N__29664));
    Span4Mux_h I__6596 (
            .O(N__29699),
            .I(N__29664));
    Span4Mux_v I__6595 (
            .O(N__29696),
            .I(N__29664));
    LocalMux I__6594 (
            .O(N__29687),
            .I(N__29664));
    Span4Mux_h I__6593 (
            .O(N__29678),
            .I(N__29661));
    Odrv4 I__6592 (
            .O(N__29673),
            .I(\this_vga_signals.GZ0Z_424 ));
    Odrv4 I__6591 (
            .O(N__29664),
            .I(\this_vga_signals.GZ0Z_424 ));
    Odrv4 I__6590 (
            .O(N__29661),
            .I(\this_vga_signals.GZ0Z_424 ));
    IoInMux I__6589 (
            .O(N__29654),
            .I(N__29651));
    LocalMux I__6588 (
            .O(N__29651),
            .I(N__29647));
    InMux I__6587 (
            .O(N__29650),
            .I(N__29644));
    Span12Mux_s8_v I__6586 (
            .O(N__29647),
            .I(N__29641));
    LocalMux I__6585 (
            .O(N__29644),
            .I(\this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9 ));
    Odrv12 I__6584 (
            .O(N__29641),
            .I(\this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9 ));
    InMux I__6583 (
            .O(N__29636),
            .I(N__29633));
    LocalMux I__6582 (
            .O(N__29633),
            .I(N__29630));
    Sp12to4 I__6581 (
            .O(N__29630),
            .I(N__29627));
    Span12Mux_v I__6580 (
            .O(N__29627),
            .I(N__29624));
    Odrv12 I__6579 (
            .O(N__29624),
            .I(\this_ppu.oam_cache.mem_1 ));
    CascadeMux I__6578 (
            .O(N__29621),
            .I(\this_vga_signals.vvisibility_0_cascade_ ));
    CascadeMux I__6577 (
            .O(N__29618),
            .I(N__29614));
    InMux I__6576 (
            .O(N__29617),
            .I(N__29611));
    InMux I__6575 (
            .O(N__29614),
            .I(N__29608));
    LocalMux I__6574 (
            .O(N__29611),
            .I(N__29602));
    LocalMux I__6573 (
            .O(N__29608),
            .I(N__29602));
    InMux I__6572 (
            .O(N__29607),
            .I(N__29599));
    Span12Mux_v I__6571 (
            .O(N__29602),
            .I(N__29595));
    LocalMux I__6570 (
            .O(N__29599),
            .I(N__29592));
    InMux I__6569 (
            .O(N__29598),
            .I(N__29589));
    Span12Mux_h I__6568 (
            .O(N__29595),
            .I(N__29586));
    Span4Mux_h I__6567 (
            .O(N__29592),
            .I(N__29583));
    LocalMux I__6566 (
            .O(N__29589),
            .I(\this_vga_signals.vvisibility ));
    Odrv12 I__6565 (
            .O(N__29586),
            .I(\this_vga_signals.vvisibility ));
    Odrv4 I__6564 (
            .O(N__29583),
            .I(\this_vga_signals.vvisibility ));
    CascadeMux I__6563 (
            .O(N__29576),
            .I(N__29566));
    CascadeMux I__6562 (
            .O(N__29575),
            .I(N__29563));
    CascadeMux I__6561 (
            .O(N__29574),
            .I(N__29559));
    CascadeMux I__6560 (
            .O(N__29573),
            .I(N__29556));
    CascadeMux I__6559 (
            .O(N__29572),
            .I(N__29552));
    CascadeMux I__6558 (
            .O(N__29571),
            .I(N__29547));
    CascadeMux I__6557 (
            .O(N__29570),
            .I(N__29543));
    CascadeMux I__6556 (
            .O(N__29569),
            .I(N__29540));
    InMux I__6555 (
            .O(N__29566),
            .I(N__29537));
    InMux I__6554 (
            .O(N__29563),
            .I(N__29534));
    CascadeMux I__6553 (
            .O(N__29562),
            .I(N__29531));
    InMux I__6552 (
            .O(N__29559),
            .I(N__29528));
    InMux I__6551 (
            .O(N__29556),
            .I(N__29525));
    CascadeMux I__6550 (
            .O(N__29555),
            .I(N__29522));
    InMux I__6549 (
            .O(N__29552),
            .I(N__29519));
    CascadeMux I__6548 (
            .O(N__29551),
            .I(N__29516));
    CascadeMux I__6547 (
            .O(N__29550),
            .I(N__29511));
    InMux I__6546 (
            .O(N__29547),
            .I(N__29508));
    CascadeMux I__6545 (
            .O(N__29546),
            .I(N__29505));
    InMux I__6544 (
            .O(N__29543),
            .I(N__29502));
    InMux I__6543 (
            .O(N__29540),
            .I(N__29499));
    LocalMux I__6542 (
            .O(N__29537),
            .I(N__29494));
    LocalMux I__6541 (
            .O(N__29534),
            .I(N__29494));
    InMux I__6540 (
            .O(N__29531),
            .I(N__29491));
    LocalMux I__6539 (
            .O(N__29528),
            .I(N__29486));
    LocalMux I__6538 (
            .O(N__29525),
            .I(N__29486));
    InMux I__6537 (
            .O(N__29522),
            .I(N__29483));
    LocalMux I__6536 (
            .O(N__29519),
            .I(N__29480));
    InMux I__6535 (
            .O(N__29516),
            .I(N__29477));
    CascadeMux I__6534 (
            .O(N__29515),
            .I(N__29474));
    CascadeMux I__6533 (
            .O(N__29514),
            .I(N__29471));
    InMux I__6532 (
            .O(N__29511),
            .I(N__29468));
    LocalMux I__6531 (
            .O(N__29508),
            .I(N__29465));
    InMux I__6530 (
            .O(N__29505),
            .I(N__29462));
    LocalMux I__6529 (
            .O(N__29502),
            .I(N__29459));
    LocalMux I__6528 (
            .O(N__29499),
            .I(N__29454));
    Span4Mux_v I__6527 (
            .O(N__29494),
            .I(N__29454));
    LocalMux I__6526 (
            .O(N__29491),
            .I(N__29449));
    Span4Mux_v I__6525 (
            .O(N__29486),
            .I(N__29449));
    LocalMux I__6524 (
            .O(N__29483),
            .I(N__29445));
    Span4Mux_v I__6523 (
            .O(N__29480),
            .I(N__29440));
    LocalMux I__6522 (
            .O(N__29477),
            .I(N__29440));
    InMux I__6521 (
            .O(N__29474),
            .I(N__29437));
    InMux I__6520 (
            .O(N__29471),
            .I(N__29434));
    LocalMux I__6519 (
            .O(N__29468),
            .I(N__29427));
    Span4Mux_s2_v I__6518 (
            .O(N__29465),
            .I(N__29427));
    LocalMux I__6517 (
            .O(N__29462),
            .I(N__29427));
    Span4Mux_v I__6516 (
            .O(N__29459),
            .I(N__29424));
    Span4Mux_v I__6515 (
            .O(N__29454),
            .I(N__29421));
    Sp12to4 I__6514 (
            .O(N__29449),
            .I(N__29418));
    CascadeMux I__6513 (
            .O(N__29448),
            .I(N__29415));
    Span4Mux_v I__6512 (
            .O(N__29445),
            .I(N__29412));
    Span4Mux_v I__6511 (
            .O(N__29440),
            .I(N__29409));
    LocalMux I__6510 (
            .O(N__29437),
            .I(N__29402));
    LocalMux I__6509 (
            .O(N__29434),
            .I(N__29402));
    Span4Mux_v I__6508 (
            .O(N__29427),
            .I(N__29402));
    Span4Mux_h I__6507 (
            .O(N__29424),
            .I(N__29396));
    Span4Mux_h I__6506 (
            .O(N__29421),
            .I(N__29396));
    Span12Mux_h I__6505 (
            .O(N__29418),
            .I(N__29393));
    InMux I__6504 (
            .O(N__29415),
            .I(N__29390));
    Sp12to4 I__6503 (
            .O(N__29412),
            .I(N__29385));
    Sp12to4 I__6502 (
            .O(N__29409),
            .I(N__29385));
    Sp12to4 I__6501 (
            .O(N__29402),
            .I(N__29382));
    InMux I__6500 (
            .O(N__29401),
            .I(N__29379));
    Span4Mux_h I__6499 (
            .O(N__29396),
            .I(N__29376));
    Span12Mux_v I__6498 (
            .O(N__29393),
            .I(N__29373));
    LocalMux I__6497 (
            .O(N__29390),
            .I(N__29366));
    Span12Mux_v I__6496 (
            .O(N__29385),
            .I(N__29366));
    Span12Mux_s11_v I__6495 (
            .O(N__29382),
            .I(N__29366));
    LocalMux I__6494 (
            .O(N__29379),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv4 I__6493 (
            .O(N__29376),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv12 I__6492 (
            .O(N__29373),
            .I(M_this_spr_address_qZ0Z_7));
    Odrv12 I__6491 (
            .O(N__29366),
            .I(M_this_spr_address_qZ0Z_7));
    InMux I__6490 (
            .O(N__29357),
            .I(un1_M_this_spr_address_q_cry_6));
    CascadeMux I__6489 (
            .O(N__29354),
            .I(N__29345));
    CascadeMux I__6488 (
            .O(N__29353),
            .I(N__29342));
    CascadeMux I__6487 (
            .O(N__29352),
            .I(N__29337));
    CascadeMux I__6486 (
            .O(N__29351),
            .I(N__29334));
    CascadeMux I__6485 (
            .O(N__29350),
            .I(N__29331));
    CascadeMux I__6484 (
            .O(N__29349),
            .I(N__29328));
    CascadeMux I__6483 (
            .O(N__29348),
            .I(N__29325));
    InMux I__6482 (
            .O(N__29345),
            .I(N__29322));
    InMux I__6481 (
            .O(N__29342),
            .I(N__29319));
    CascadeMux I__6480 (
            .O(N__29341),
            .I(N__29315));
    CascadeMux I__6479 (
            .O(N__29340),
            .I(N__29312));
    InMux I__6478 (
            .O(N__29337),
            .I(N__29308));
    InMux I__6477 (
            .O(N__29334),
            .I(N__29305));
    InMux I__6476 (
            .O(N__29331),
            .I(N__29302));
    InMux I__6475 (
            .O(N__29328),
            .I(N__29299));
    InMux I__6474 (
            .O(N__29325),
            .I(N__29296));
    LocalMux I__6473 (
            .O(N__29322),
            .I(N__29293));
    LocalMux I__6472 (
            .O(N__29319),
            .I(N__29290));
    CascadeMux I__6471 (
            .O(N__29318),
            .I(N__29282));
    InMux I__6470 (
            .O(N__29315),
            .I(N__29279));
    InMux I__6469 (
            .O(N__29312),
            .I(N__29276));
    CascadeMux I__6468 (
            .O(N__29311),
            .I(N__29273));
    LocalMux I__6467 (
            .O(N__29308),
            .I(N__29268));
    LocalMux I__6466 (
            .O(N__29305),
            .I(N__29268));
    LocalMux I__6465 (
            .O(N__29302),
            .I(N__29265));
    LocalMux I__6464 (
            .O(N__29299),
            .I(N__29260));
    LocalMux I__6463 (
            .O(N__29296),
            .I(N__29260));
    Span4Mux_v I__6462 (
            .O(N__29293),
            .I(N__29255));
    Span4Mux_v I__6461 (
            .O(N__29290),
            .I(N__29255));
    CascadeMux I__6460 (
            .O(N__29289),
            .I(N__29252));
    CascadeMux I__6459 (
            .O(N__29288),
            .I(N__29249));
    CascadeMux I__6458 (
            .O(N__29287),
            .I(N__29246));
    CascadeMux I__6457 (
            .O(N__29286),
            .I(N__29243));
    CascadeMux I__6456 (
            .O(N__29285),
            .I(N__29240));
    InMux I__6455 (
            .O(N__29282),
            .I(N__29237));
    LocalMux I__6454 (
            .O(N__29279),
            .I(N__29232));
    LocalMux I__6453 (
            .O(N__29276),
            .I(N__29232));
    InMux I__6452 (
            .O(N__29273),
            .I(N__29229));
    Span4Mux_v I__6451 (
            .O(N__29268),
            .I(N__29224));
    Span4Mux_v I__6450 (
            .O(N__29265),
            .I(N__29224));
    Span4Mux_v I__6449 (
            .O(N__29260),
            .I(N__29221));
    Span4Mux_v I__6448 (
            .O(N__29255),
            .I(N__29218));
    InMux I__6447 (
            .O(N__29252),
            .I(N__29215));
    InMux I__6446 (
            .O(N__29249),
            .I(N__29212));
    InMux I__6445 (
            .O(N__29246),
            .I(N__29209));
    InMux I__6444 (
            .O(N__29243),
            .I(N__29206));
    InMux I__6443 (
            .O(N__29240),
            .I(N__29203));
    LocalMux I__6442 (
            .O(N__29237),
            .I(N__29196));
    Span4Mux_v I__6441 (
            .O(N__29232),
            .I(N__29196));
    LocalMux I__6440 (
            .O(N__29229),
            .I(N__29196));
    Span4Mux_h I__6439 (
            .O(N__29224),
            .I(N__29193));
    Span4Mux_h I__6438 (
            .O(N__29221),
            .I(N__29187));
    Span4Mux_h I__6437 (
            .O(N__29218),
            .I(N__29187));
    LocalMux I__6436 (
            .O(N__29215),
            .I(N__29180));
    LocalMux I__6435 (
            .O(N__29212),
            .I(N__29180));
    LocalMux I__6434 (
            .O(N__29209),
            .I(N__29180));
    LocalMux I__6433 (
            .O(N__29206),
            .I(N__29173));
    LocalMux I__6432 (
            .O(N__29203),
            .I(N__29173));
    Sp12to4 I__6431 (
            .O(N__29196),
            .I(N__29173));
    Sp12to4 I__6430 (
            .O(N__29193),
            .I(N__29170));
    InMux I__6429 (
            .O(N__29192),
            .I(N__29167));
    Span4Mux_h I__6428 (
            .O(N__29187),
            .I(N__29164));
    Span12Mux_v I__6427 (
            .O(N__29180),
            .I(N__29157));
    Span12Mux_v I__6426 (
            .O(N__29173),
            .I(N__29157));
    Span12Mux_v I__6425 (
            .O(N__29170),
            .I(N__29157));
    LocalMux I__6424 (
            .O(N__29167),
            .I(M_this_spr_address_qZ0Z_8));
    Odrv4 I__6423 (
            .O(N__29164),
            .I(M_this_spr_address_qZ0Z_8));
    Odrv12 I__6422 (
            .O(N__29157),
            .I(M_this_spr_address_qZ0Z_8));
    InMux I__6421 (
            .O(N__29150),
            .I(bfn_17_13_0_));
    CascadeMux I__6420 (
            .O(N__29147),
            .I(N__29144));
    InMux I__6419 (
            .O(N__29144),
            .I(N__29139));
    CascadeMux I__6418 (
            .O(N__29143),
            .I(N__29136));
    CascadeMux I__6417 (
            .O(N__29142),
            .I(N__29132));
    LocalMux I__6416 (
            .O(N__29139),
            .I(N__29129));
    InMux I__6415 (
            .O(N__29136),
            .I(N__29126));
    CascadeMux I__6414 (
            .O(N__29135),
            .I(N__29123));
    InMux I__6413 (
            .O(N__29132),
            .I(N__29117));
    Span4Mux_h I__6412 (
            .O(N__29129),
            .I(N__29112));
    LocalMux I__6411 (
            .O(N__29126),
            .I(N__29112));
    InMux I__6410 (
            .O(N__29123),
            .I(N__29109));
    CascadeMux I__6409 (
            .O(N__29122),
            .I(N__29106));
    CascadeMux I__6408 (
            .O(N__29121),
            .I(N__29102));
    CascadeMux I__6407 (
            .O(N__29120),
            .I(N__29095));
    LocalMux I__6406 (
            .O(N__29117),
            .I(N__29088));
    Span4Mux_v I__6405 (
            .O(N__29112),
            .I(N__29088));
    LocalMux I__6404 (
            .O(N__29109),
            .I(N__29088));
    InMux I__6403 (
            .O(N__29106),
            .I(N__29085));
    CascadeMux I__6402 (
            .O(N__29105),
            .I(N__29082));
    InMux I__6401 (
            .O(N__29102),
            .I(N__29077));
    CascadeMux I__6400 (
            .O(N__29101),
            .I(N__29074));
    CascadeMux I__6399 (
            .O(N__29100),
            .I(N__29071));
    CascadeMux I__6398 (
            .O(N__29099),
            .I(N__29068));
    CascadeMux I__6397 (
            .O(N__29098),
            .I(N__29065));
    InMux I__6396 (
            .O(N__29095),
            .I(N__29062));
    Span4Mux_v I__6395 (
            .O(N__29088),
            .I(N__29057));
    LocalMux I__6394 (
            .O(N__29085),
            .I(N__29057));
    InMux I__6393 (
            .O(N__29082),
            .I(N__29054));
    CascadeMux I__6392 (
            .O(N__29081),
            .I(N__29051));
    CascadeMux I__6391 (
            .O(N__29080),
            .I(N__29048));
    LocalMux I__6390 (
            .O(N__29077),
            .I(N__29044));
    InMux I__6389 (
            .O(N__29074),
            .I(N__29041));
    InMux I__6388 (
            .O(N__29071),
            .I(N__29038));
    InMux I__6387 (
            .O(N__29068),
            .I(N__29035));
    InMux I__6386 (
            .O(N__29065),
            .I(N__29032));
    LocalMux I__6385 (
            .O(N__29062),
            .I(N__29029));
    Span4Mux_h I__6384 (
            .O(N__29057),
            .I(N__29023));
    LocalMux I__6383 (
            .O(N__29054),
            .I(N__29023));
    InMux I__6382 (
            .O(N__29051),
            .I(N__29020));
    InMux I__6381 (
            .O(N__29048),
            .I(N__29017));
    CascadeMux I__6380 (
            .O(N__29047),
            .I(N__29014));
    Span4Mux_v I__6379 (
            .O(N__29044),
            .I(N__29011));
    LocalMux I__6378 (
            .O(N__29041),
            .I(N__29006));
    LocalMux I__6377 (
            .O(N__29038),
            .I(N__29006));
    LocalMux I__6376 (
            .O(N__29035),
            .I(N__29003));
    LocalMux I__6375 (
            .O(N__29032),
            .I(N__29000));
    Span4Mux_h I__6374 (
            .O(N__29029),
            .I(N__28997));
    CascadeMux I__6373 (
            .O(N__29028),
            .I(N__28994));
    Span4Mux_v I__6372 (
            .O(N__29023),
            .I(N__28987));
    LocalMux I__6371 (
            .O(N__29020),
            .I(N__28987));
    LocalMux I__6370 (
            .O(N__29017),
            .I(N__28987));
    InMux I__6369 (
            .O(N__29014),
            .I(N__28984));
    Span4Mux_h I__6368 (
            .O(N__29011),
            .I(N__28981));
    Span4Mux_v I__6367 (
            .O(N__29006),
            .I(N__28978));
    Span4Mux_h I__6366 (
            .O(N__29003),
            .I(N__28975));
    Span4Mux_h I__6365 (
            .O(N__29000),
            .I(N__28972));
    Sp12to4 I__6364 (
            .O(N__28997),
            .I(N__28969));
    InMux I__6363 (
            .O(N__28994),
            .I(N__28966));
    Span4Mux_v I__6362 (
            .O(N__28987),
            .I(N__28963));
    LocalMux I__6361 (
            .O(N__28984),
            .I(N__28960));
    Span4Mux_v I__6360 (
            .O(N__28981),
            .I(N__28954));
    Span4Mux_h I__6359 (
            .O(N__28978),
            .I(N__28954));
    Sp12to4 I__6358 (
            .O(N__28975),
            .I(N__28947));
    Sp12to4 I__6357 (
            .O(N__28972),
            .I(N__28947));
    Span12Mux_s7_v I__6356 (
            .O(N__28969),
            .I(N__28947));
    LocalMux I__6355 (
            .O(N__28966),
            .I(N__28944));
    Sp12to4 I__6354 (
            .O(N__28963),
            .I(N__28939));
    Sp12to4 I__6353 (
            .O(N__28960),
            .I(N__28939));
    InMux I__6352 (
            .O(N__28959),
            .I(N__28936));
    Span4Mux_h I__6351 (
            .O(N__28954),
            .I(N__28933));
    Span12Mux_v I__6350 (
            .O(N__28947),
            .I(N__28930));
    Span12Mux_h I__6349 (
            .O(N__28944),
            .I(N__28925));
    Span12Mux_h I__6348 (
            .O(N__28939),
            .I(N__28925));
    LocalMux I__6347 (
            .O(N__28936),
            .I(M_this_spr_address_qZ0Z_9));
    Odrv4 I__6346 (
            .O(N__28933),
            .I(M_this_spr_address_qZ0Z_9));
    Odrv12 I__6345 (
            .O(N__28930),
            .I(M_this_spr_address_qZ0Z_9));
    Odrv12 I__6344 (
            .O(N__28925),
            .I(M_this_spr_address_qZ0Z_9));
    InMux I__6343 (
            .O(N__28916),
            .I(un1_M_this_spr_address_q_cry_8));
    CascadeMux I__6342 (
            .O(N__28913),
            .I(N__28908));
    CascadeMux I__6341 (
            .O(N__28912),
            .I(N__28904));
    CascadeMux I__6340 (
            .O(N__28911),
            .I(N__28895));
    InMux I__6339 (
            .O(N__28908),
            .I(N__28891));
    CascadeMux I__6338 (
            .O(N__28907),
            .I(N__28887));
    InMux I__6337 (
            .O(N__28904),
            .I(N__28884));
    CascadeMux I__6336 (
            .O(N__28903),
            .I(N__28881));
    CascadeMux I__6335 (
            .O(N__28902),
            .I(N__28878));
    CascadeMux I__6334 (
            .O(N__28901),
            .I(N__28874));
    CascadeMux I__6333 (
            .O(N__28900),
            .I(N__28871));
    CascadeMux I__6332 (
            .O(N__28899),
            .I(N__28865));
    CascadeMux I__6331 (
            .O(N__28898),
            .I(N__28862));
    InMux I__6330 (
            .O(N__28895),
            .I(N__28859));
    CascadeMux I__6329 (
            .O(N__28894),
            .I(N__28856));
    LocalMux I__6328 (
            .O(N__28891),
            .I(N__28853));
    CascadeMux I__6327 (
            .O(N__28890),
            .I(N__28850));
    InMux I__6326 (
            .O(N__28887),
            .I(N__28847));
    LocalMux I__6325 (
            .O(N__28884),
            .I(N__28844));
    InMux I__6324 (
            .O(N__28881),
            .I(N__28841));
    InMux I__6323 (
            .O(N__28878),
            .I(N__28838));
    CascadeMux I__6322 (
            .O(N__28877),
            .I(N__28835));
    InMux I__6321 (
            .O(N__28874),
            .I(N__28832));
    InMux I__6320 (
            .O(N__28871),
            .I(N__28829));
    CascadeMux I__6319 (
            .O(N__28870),
            .I(N__28826));
    CascadeMux I__6318 (
            .O(N__28869),
            .I(N__28823));
    CascadeMux I__6317 (
            .O(N__28868),
            .I(N__28820));
    InMux I__6316 (
            .O(N__28865),
            .I(N__28817));
    InMux I__6315 (
            .O(N__28862),
            .I(N__28814));
    LocalMux I__6314 (
            .O(N__28859),
            .I(N__28811));
    InMux I__6313 (
            .O(N__28856),
            .I(N__28808));
    Span4Mux_v I__6312 (
            .O(N__28853),
            .I(N__28805));
    InMux I__6311 (
            .O(N__28850),
            .I(N__28802));
    LocalMux I__6310 (
            .O(N__28847),
            .I(N__28799));
    Span4Mux_v I__6309 (
            .O(N__28844),
            .I(N__28792));
    LocalMux I__6308 (
            .O(N__28841),
            .I(N__28792));
    LocalMux I__6307 (
            .O(N__28838),
            .I(N__28792));
    InMux I__6306 (
            .O(N__28835),
            .I(N__28789));
    LocalMux I__6305 (
            .O(N__28832),
            .I(N__28784));
    LocalMux I__6304 (
            .O(N__28829),
            .I(N__28784));
    InMux I__6303 (
            .O(N__28826),
            .I(N__28781));
    InMux I__6302 (
            .O(N__28823),
            .I(N__28778));
    InMux I__6301 (
            .O(N__28820),
            .I(N__28775));
    LocalMux I__6300 (
            .O(N__28817),
            .I(N__28772));
    LocalMux I__6299 (
            .O(N__28814),
            .I(N__28767));
    Span4Mux_h I__6298 (
            .O(N__28811),
            .I(N__28767));
    LocalMux I__6297 (
            .O(N__28808),
            .I(N__28764));
    Span4Mux_h I__6296 (
            .O(N__28805),
            .I(N__28757));
    LocalMux I__6295 (
            .O(N__28802),
            .I(N__28757));
    Span4Mux_v I__6294 (
            .O(N__28799),
            .I(N__28757));
    Span4Mux_v I__6293 (
            .O(N__28792),
            .I(N__28752));
    LocalMux I__6292 (
            .O(N__28789),
            .I(N__28752));
    Span4Mux_v I__6291 (
            .O(N__28784),
            .I(N__28745));
    LocalMux I__6290 (
            .O(N__28781),
            .I(N__28745));
    LocalMux I__6289 (
            .O(N__28778),
            .I(N__28745));
    LocalMux I__6288 (
            .O(N__28775),
            .I(N__28742));
    Span4Mux_h I__6287 (
            .O(N__28772),
            .I(N__28735));
    Span4Mux_v I__6286 (
            .O(N__28767),
            .I(N__28735));
    Span4Mux_v I__6285 (
            .O(N__28764),
            .I(N__28735));
    Span4Mux_v I__6284 (
            .O(N__28757),
            .I(N__28732));
    Span4Mux_s2_v I__6283 (
            .O(N__28752),
            .I(N__28729));
    Span4Mux_v I__6282 (
            .O(N__28745),
            .I(N__28726));
    Span4Mux_s2_v I__6281 (
            .O(N__28742),
            .I(N__28723));
    Span4Mux_h I__6280 (
            .O(N__28735),
            .I(N__28719));
    Sp12to4 I__6279 (
            .O(N__28732),
            .I(N__28716));
    Sp12to4 I__6278 (
            .O(N__28729),
            .I(N__28713));
    Sp12to4 I__6277 (
            .O(N__28726),
            .I(N__28708));
    Sp12to4 I__6276 (
            .O(N__28723),
            .I(N__28708));
    InMux I__6275 (
            .O(N__28722),
            .I(N__28705));
    Span4Mux_h I__6274 (
            .O(N__28719),
            .I(N__28702));
    Span12Mux_h I__6273 (
            .O(N__28716),
            .I(N__28699));
    Span12Mux_h I__6272 (
            .O(N__28713),
            .I(N__28694));
    Span12Mux_h I__6271 (
            .O(N__28708),
            .I(N__28694));
    LocalMux I__6270 (
            .O(N__28705),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv4 I__6269 (
            .O(N__28702),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv12 I__6268 (
            .O(N__28699),
            .I(M_this_spr_address_qZ0Z_10));
    Odrv12 I__6267 (
            .O(N__28694),
            .I(M_this_spr_address_qZ0Z_10));
    InMux I__6266 (
            .O(N__28685),
            .I(un1_M_this_spr_address_q_cry_9));
    InMux I__6265 (
            .O(N__28682),
            .I(un1_M_this_spr_address_q_cry_10));
    InMux I__6264 (
            .O(N__28679),
            .I(un1_M_this_spr_address_q_cry_11));
    InMux I__6263 (
            .O(N__28676),
            .I(un1_M_this_spr_address_q_cry_12));
    CascadeMux I__6262 (
            .O(N__28673),
            .I(N__28669));
    InMux I__6261 (
            .O(N__28672),
            .I(N__28666));
    InMux I__6260 (
            .O(N__28669),
            .I(N__28663));
    LocalMux I__6259 (
            .O(N__28666),
            .I(N__28658));
    LocalMux I__6258 (
            .O(N__28663),
            .I(N__28658));
    Odrv4 I__6257 (
            .O(N__28658),
            .I(M_this_spr_ram_write_en_0_i_1));
    InMux I__6256 (
            .O(N__28655),
            .I(N__28651));
    InMux I__6255 (
            .O(N__28654),
            .I(N__28648));
    LocalMux I__6254 (
            .O(N__28651),
            .I(N__28644));
    LocalMux I__6253 (
            .O(N__28648),
            .I(N__28641));
    InMux I__6252 (
            .O(N__28647),
            .I(N__28638));
    Span4Mux_v I__6251 (
            .O(N__28644),
            .I(N__28635));
    Span4Mux_v I__6250 (
            .O(N__28641),
            .I(N__28632));
    LocalMux I__6249 (
            .O(N__28638),
            .I(N__28629));
    Span4Mux_h I__6248 (
            .O(N__28635),
            .I(N__28626));
    Span4Mux_h I__6247 (
            .O(N__28632),
            .I(N__28621));
    Span4Mux_h I__6246 (
            .O(N__28629),
            .I(N__28621));
    Odrv4 I__6245 (
            .O(N__28626),
            .I(\this_vga_signals.M_vcounter_d8 ));
    Odrv4 I__6244 (
            .O(N__28621),
            .I(\this_vga_signals.M_vcounter_d8 ));
    CascadeMux I__6243 (
            .O(N__28616),
            .I(N__28607));
    InMux I__6242 (
            .O(N__28615),
            .I(N__28604));
    InMux I__6241 (
            .O(N__28614),
            .I(N__28597));
    InMux I__6240 (
            .O(N__28613),
            .I(N__28597));
    InMux I__6239 (
            .O(N__28612),
            .I(N__28597));
    InMux I__6238 (
            .O(N__28611),
            .I(N__28593));
    InMux I__6237 (
            .O(N__28610),
            .I(N__28590));
    InMux I__6236 (
            .O(N__28607),
            .I(N__28587));
    LocalMux I__6235 (
            .O(N__28604),
            .I(N__28583));
    LocalMux I__6234 (
            .O(N__28597),
            .I(N__28580));
    InMux I__6233 (
            .O(N__28596),
            .I(N__28577));
    LocalMux I__6232 (
            .O(N__28593),
            .I(N__28570));
    LocalMux I__6231 (
            .O(N__28590),
            .I(N__28570));
    LocalMux I__6230 (
            .O(N__28587),
            .I(N__28570));
    InMux I__6229 (
            .O(N__28586),
            .I(N__28564));
    Span4Mux_v I__6228 (
            .O(N__28583),
            .I(N__28557));
    Span4Mux_h I__6227 (
            .O(N__28580),
            .I(N__28557));
    LocalMux I__6226 (
            .O(N__28577),
            .I(N__28557));
    Span12Mux_h I__6225 (
            .O(N__28570),
            .I(N__28554));
    InMux I__6224 (
            .O(N__28569),
            .I(N__28547));
    InMux I__6223 (
            .O(N__28568),
            .I(N__28547));
    InMux I__6222 (
            .O(N__28567),
            .I(N__28547));
    LocalMux I__6221 (
            .O(N__28564),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv4 I__6220 (
            .O(N__28557),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    Odrv12 I__6219 (
            .O(N__28554),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    LocalMux I__6218 (
            .O(N__28547),
            .I(\this_vga_signals.M_hcounter_d7_0 ));
    InMux I__6217 (
            .O(N__28538),
            .I(N__28535));
    LocalMux I__6216 (
            .O(N__28535),
            .I(N__28531));
    CascadeMux I__6215 (
            .O(N__28534),
            .I(N__28528));
    Span4Mux_v I__6214 (
            .O(N__28531),
            .I(N__28525));
    InMux I__6213 (
            .O(N__28528),
            .I(N__28522));
    Odrv4 I__6212 (
            .O(N__28525),
            .I(M_this_ctrl_flags_qZ0Z_7));
    LocalMux I__6211 (
            .O(N__28522),
            .I(M_this_ctrl_flags_qZ0Z_7));
    InMux I__6210 (
            .O(N__28517),
            .I(N__28514));
    LocalMux I__6209 (
            .O(N__28514),
            .I(N__28511));
    Odrv4 I__6208 (
            .O(N__28511),
            .I(\this_reset_cond.M_stage_qZ0Z_5 ));
    CascadeMux I__6207 (
            .O(N__28508),
            .I(N__28502));
    CascadeMux I__6206 (
            .O(N__28507),
            .I(N__28499));
    CascadeMux I__6205 (
            .O(N__28506),
            .I(N__28496));
    CascadeMux I__6204 (
            .O(N__28505),
            .I(N__28492));
    InMux I__6203 (
            .O(N__28502),
            .I(N__28487));
    InMux I__6202 (
            .O(N__28499),
            .I(N__28484));
    InMux I__6201 (
            .O(N__28496),
            .I(N__28481));
    CascadeMux I__6200 (
            .O(N__28495),
            .I(N__28478));
    InMux I__6199 (
            .O(N__28492),
            .I(N__28474));
    CascadeMux I__6198 (
            .O(N__28491),
            .I(N__28471));
    CascadeMux I__6197 (
            .O(N__28490),
            .I(N__28466));
    LocalMux I__6196 (
            .O(N__28487),
            .I(N__28460));
    LocalMux I__6195 (
            .O(N__28484),
            .I(N__28460));
    LocalMux I__6194 (
            .O(N__28481),
            .I(N__28456));
    InMux I__6193 (
            .O(N__28478),
            .I(N__28453));
    CascadeMux I__6192 (
            .O(N__28477),
            .I(N__28450));
    LocalMux I__6191 (
            .O(N__28474),
            .I(N__28447));
    InMux I__6190 (
            .O(N__28471),
            .I(N__28444));
    CascadeMux I__6189 (
            .O(N__28470),
            .I(N__28441));
    CascadeMux I__6188 (
            .O(N__28469),
            .I(N__28438));
    InMux I__6187 (
            .O(N__28466),
            .I(N__28434));
    CascadeMux I__6186 (
            .O(N__28465),
            .I(N__28431));
    Span4Mux_v I__6185 (
            .O(N__28460),
            .I(N__28426));
    CascadeMux I__6184 (
            .O(N__28459),
            .I(N__28423));
    Span4Mux_s3_v I__6183 (
            .O(N__28456),
            .I(N__28418));
    LocalMux I__6182 (
            .O(N__28453),
            .I(N__28418));
    InMux I__6181 (
            .O(N__28450),
            .I(N__28415));
    Span4Mux_s1_v I__6180 (
            .O(N__28447),
            .I(N__28409));
    LocalMux I__6179 (
            .O(N__28444),
            .I(N__28409));
    InMux I__6178 (
            .O(N__28441),
            .I(N__28406));
    InMux I__6177 (
            .O(N__28438),
            .I(N__28403));
    CascadeMux I__6176 (
            .O(N__28437),
            .I(N__28400));
    LocalMux I__6175 (
            .O(N__28434),
            .I(N__28397));
    InMux I__6174 (
            .O(N__28431),
            .I(N__28394));
    CascadeMux I__6173 (
            .O(N__28430),
            .I(N__28391));
    CascadeMux I__6172 (
            .O(N__28429),
            .I(N__28388));
    Span4Mux_h I__6171 (
            .O(N__28426),
            .I(N__28385));
    InMux I__6170 (
            .O(N__28423),
            .I(N__28382));
    Span4Mux_h I__6169 (
            .O(N__28418),
            .I(N__28377));
    LocalMux I__6168 (
            .O(N__28415),
            .I(N__28377));
    CascadeMux I__6167 (
            .O(N__28414),
            .I(N__28374));
    Span4Mux_v I__6166 (
            .O(N__28409),
            .I(N__28369));
    LocalMux I__6165 (
            .O(N__28406),
            .I(N__28369));
    LocalMux I__6164 (
            .O(N__28403),
            .I(N__28366));
    InMux I__6163 (
            .O(N__28400),
            .I(N__28363));
    Span4Mux_h I__6162 (
            .O(N__28397),
            .I(N__28358));
    LocalMux I__6161 (
            .O(N__28394),
            .I(N__28358));
    InMux I__6160 (
            .O(N__28391),
            .I(N__28355));
    InMux I__6159 (
            .O(N__28388),
            .I(N__28352));
    Span4Mux_h I__6158 (
            .O(N__28385),
            .I(N__28349));
    LocalMux I__6157 (
            .O(N__28382),
            .I(N__28346));
    Span4Mux_v I__6156 (
            .O(N__28377),
            .I(N__28343));
    InMux I__6155 (
            .O(N__28374),
            .I(N__28340));
    Span4Mux_h I__6154 (
            .O(N__28369),
            .I(N__28337));
    Span4Mux_v I__6153 (
            .O(N__28366),
            .I(N__28332));
    LocalMux I__6152 (
            .O(N__28363),
            .I(N__28332));
    Span4Mux_v I__6151 (
            .O(N__28358),
            .I(N__28327));
    LocalMux I__6150 (
            .O(N__28355),
            .I(N__28327));
    LocalMux I__6149 (
            .O(N__28352),
            .I(N__28324));
    Sp12to4 I__6148 (
            .O(N__28349),
            .I(N__28319));
    Span12Mux_h I__6147 (
            .O(N__28346),
            .I(N__28319));
    Sp12to4 I__6146 (
            .O(N__28343),
            .I(N__28314));
    LocalMux I__6145 (
            .O(N__28340),
            .I(N__28314));
    Span4Mux_v I__6144 (
            .O(N__28337),
            .I(N__28309));
    Span4Mux_h I__6143 (
            .O(N__28332),
            .I(N__28309));
    Span4Mux_h I__6142 (
            .O(N__28327),
            .I(N__28306));
    Span4Mux_h I__6141 (
            .O(N__28324),
            .I(N__28303));
    Span12Mux_v I__6140 (
            .O(N__28319),
            .I(N__28299));
    Span12Mux_h I__6139 (
            .O(N__28314),
            .I(N__28296));
    Span4Mux_h I__6138 (
            .O(N__28309),
            .I(N__28291));
    Span4Mux_h I__6137 (
            .O(N__28306),
            .I(N__28291));
    Span4Mux_h I__6136 (
            .O(N__28303),
            .I(N__28288));
    InMux I__6135 (
            .O(N__28302),
            .I(N__28285));
    Odrv12 I__6134 (
            .O(N__28299),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv12 I__6133 (
            .O(N__28296),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv4 I__6132 (
            .O(N__28291),
            .I(M_this_spr_address_qZ0Z_0));
    Odrv4 I__6131 (
            .O(N__28288),
            .I(M_this_spr_address_qZ0Z_0));
    LocalMux I__6130 (
            .O(N__28285),
            .I(M_this_spr_address_qZ0Z_0));
    CascadeMux I__6129 (
            .O(N__28274),
            .I(N__28271));
    InMux I__6128 (
            .O(N__28271),
            .I(N__28266));
    CascadeMux I__6127 (
            .O(N__28270),
            .I(N__28263));
    CascadeMux I__6126 (
            .O(N__28269),
            .I(N__28258));
    LocalMux I__6125 (
            .O(N__28266),
            .I(N__28254));
    InMux I__6124 (
            .O(N__28263),
            .I(N__28251));
    CascadeMux I__6123 (
            .O(N__28262),
            .I(N__28248));
    CascadeMux I__6122 (
            .O(N__28261),
            .I(N__28244));
    InMux I__6121 (
            .O(N__28258),
            .I(N__28240));
    CascadeMux I__6120 (
            .O(N__28257),
            .I(N__28237));
    Span4Mux_s3_v I__6119 (
            .O(N__28254),
            .I(N__28230));
    LocalMux I__6118 (
            .O(N__28251),
            .I(N__28230));
    InMux I__6117 (
            .O(N__28248),
            .I(N__28227));
    CascadeMux I__6116 (
            .O(N__28247),
            .I(N__28224));
    InMux I__6115 (
            .O(N__28244),
            .I(N__28220));
    CascadeMux I__6114 (
            .O(N__28243),
            .I(N__28217));
    LocalMux I__6113 (
            .O(N__28240),
            .I(N__28214));
    InMux I__6112 (
            .O(N__28237),
            .I(N__28211));
    CascadeMux I__6111 (
            .O(N__28236),
            .I(N__28208));
    CascadeMux I__6110 (
            .O(N__28235),
            .I(N__28204));
    Span4Mux_h I__6109 (
            .O(N__28230),
            .I(N__28198));
    LocalMux I__6108 (
            .O(N__28227),
            .I(N__28198));
    InMux I__6107 (
            .O(N__28224),
            .I(N__28195));
    CascadeMux I__6106 (
            .O(N__28223),
            .I(N__28192));
    LocalMux I__6105 (
            .O(N__28220),
            .I(N__28188));
    InMux I__6104 (
            .O(N__28217),
            .I(N__28185));
    Span4Mux_s3_v I__6103 (
            .O(N__28214),
            .I(N__28179));
    LocalMux I__6102 (
            .O(N__28211),
            .I(N__28179));
    InMux I__6101 (
            .O(N__28208),
            .I(N__28176));
    CascadeMux I__6100 (
            .O(N__28207),
            .I(N__28173));
    InMux I__6099 (
            .O(N__28204),
            .I(N__28170));
    CascadeMux I__6098 (
            .O(N__28203),
            .I(N__28167));
    Span4Mux_v I__6097 (
            .O(N__28198),
            .I(N__28162));
    LocalMux I__6096 (
            .O(N__28195),
            .I(N__28162));
    InMux I__6095 (
            .O(N__28192),
            .I(N__28159));
    CascadeMux I__6094 (
            .O(N__28191),
            .I(N__28156));
    Span4Mux_v I__6093 (
            .O(N__28188),
            .I(N__28151));
    LocalMux I__6092 (
            .O(N__28185),
            .I(N__28151));
    CascadeMux I__6091 (
            .O(N__28184),
            .I(N__28148));
    Span4Mux_h I__6090 (
            .O(N__28179),
            .I(N__28143));
    LocalMux I__6089 (
            .O(N__28176),
            .I(N__28143));
    InMux I__6088 (
            .O(N__28173),
            .I(N__28140));
    LocalMux I__6087 (
            .O(N__28170),
            .I(N__28137));
    InMux I__6086 (
            .O(N__28167),
            .I(N__28134));
    Span4Mux_h I__6085 (
            .O(N__28162),
            .I(N__28129));
    LocalMux I__6084 (
            .O(N__28159),
            .I(N__28129));
    InMux I__6083 (
            .O(N__28156),
            .I(N__28126));
    Span4Mux_v I__6082 (
            .O(N__28151),
            .I(N__28122));
    InMux I__6081 (
            .O(N__28148),
            .I(N__28119));
    Span4Mux_v I__6080 (
            .O(N__28143),
            .I(N__28114));
    LocalMux I__6079 (
            .O(N__28140),
            .I(N__28114));
    Span4Mux_v I__6078 (
            .O(N__28137),
            .I(N__28105));
    LocalMux I__6077 (
            .O(N__28134),
            .I(N__28105));
    Span4Mux_v I__6076 (
            .O(N__28129),
            .I(N__28105));
    LocalMux I__6075 (
            .O(N__28126),
            .I(N__28105));
    CascadeMux I__6074 (
            .O(N__28125),
            .I(N__28102));
    Span4Mux_h I__6073 (
            .O(N__28122),
            .I(N__28099));
    LocalMux I__6072 (
            .O(N__28119),
            .I(N__28096));
    Span4Mux_h I__6071 (
            .O(N__28114),
            .I(N__28093));
    Span4Mux_v I__6070 (
            .O(N__28105),
            .I(N__28090));
    InMux I__6069 (
            .O(N__28102),
            .I(N__28087));
    Sp12to4 I__6068 (
            .O(N__28099),
            .I(N__28082));
    Span12Mux_s11_h I__6067 (
            .O(N__28096),
            .I(N__28082));
    Span4Mux_v I__6066 (
            .O(N__28093),
            .I(N__28079));
    Sp12to4 I__6065 (
            .O(N__28090),
            .I(N__28074));
    LocalMux I__6064 (
            .O(N__28087),
            .I(N__28074));
    Span12Mux_v I__6063 (
            .O(N__28082),
            .I(N__28066));
    Sp12to4 I__6062 (
            .O(N__28079),
            .I(N__28066));
    Span12Mux_s8_h I__6061 (
            .O(N__28074),
            .I(N__28066));
    InMux I__6060 (
            .O(N__28073),
            .I(N__28063));
    Odrv12 I__6059 (
            .O(N__28066),
            .I(M_this_spr_address_qZ0Z_1));
    LocalMux I__6058 (
            .O(N__28063),
            .I(M_this_spr_address_qZ0Z_1));
    InMux I__6057 (
            .O(N__28058),
            .I(un1_M_this_spr_address_q_cry_0));
    CascadeMux I__6056 (
            .O(N__28055),
            .I(N__28045));
    CascadeMux I__6055 (
            .O(N__28054),
            .I(N__28042));
    CascadeMux I__6054 (
            .O(N__28053),
            .I(N__28038));
    CascadeMux I__6053 (
            .O(N__28052),
            .I(N__28033));
    CascadeMux I__6052 (
            .O(N__28051),
            .I(N__28028));
    CascadeMux I__6051 (
            .O(N__28050),
            .I(N__28025));
    CascadeMux I__6050 (
            .O(N__28049),
            .I(N__28022));
    CascadeMux I__6049 (
            .O(N__28048),
            .I(N__28019));
    InMux I__6048 (
            .O(N__28045),
            .I(N__28016));
    InMux I__6047 (
            .O(N__28042),
            .I(N__28013));
    CascadeMux I__6046 (
            .O(N__28041),
            .I(N__28010));
    InMux I__6045 (
            .O(N__28038),
            .I(N__28007));
    CascadeMux I__6044 (
            .O(N__28037),
            .I(N__28001));
    CascadeMux I__6043 (
            .O(N__28036),
            .I(N__27998));
    InMux I__6042 (
            .O(N__28033),
            .I(N__27995));
    CascadeMux I__6041 (
            .O(N__28032),
            .I(N__27992));
    CascadeMux I__6040 (
            .O(N__28031),
            .I(N__27989));
    InMux I__6039 (
            .O(N__28028),
            .I(N__27986));
    InMux I__6038 (
            .O(N__28025),
            .I(N__27983));
    InMux I__6037 (
            .O(N__28022),
            .I(N__27980));
    InMux I__6036 (
            .O(N__28019),
            .I(N__27977));
    LocalMux I__6035 (
            .O(N__28016),
            .I(N__27974));
    LocalMux I__6034 (
            .O(N__28013),
            .I(N__27971));
    InMux I__6033 (
            .O(N__28010),
            .I(N__27968));
    LocalMux I__6032 (
            .O(N__28007),
            .I(N__27965));
    CascadeMux I__6031 (
            .O(N__28006),
            .I(N__27962));
    CascadeMux I__6030 (
            .O(N__28005),
            .I(N__27959));
    CascadeMux I__6029 (
            .O(N__28004),
            .I(N__27956));
    InMux I__6028 (
            .O(N__28001),
            .I(N__27953));
    InMux I__6027 (
            .O(N__27998),
            .I(N__27950));
    LocalMux I__6026 (
            .O(N__27995),
            .I(N__27947));
    InMux I__6025 (
            .O(N__27992),
            .I(N__27944));
    InMux I__6024 (
            .O(N__27989),
            .I(N__27941));
    LocalMux I__6023 (
            .O(N__27986),
            .I(N__27938));
    LocalMux I__6022 (
            .O(N__27983),
            .I(N__27935));
    LocalMux I__6021 (
            .O(N__27980),
            .I(N__27932));
    LocalMux I__6020 (
            .O(N__27977),
            .I(N__27929));
    Span4Mux_h I__6019 (
            .O(N__27974),
            .I(N__27926));
    Span4Mux_h I__6018 (
            .O(N__27971),
            .I(N__27923));
    LocalMux I__6017 (
            .O(N__27968),
            .I(N__27920));
    Span4Mux_h I__6016 (
            .O(N__27965),
            .I(N__27917));
    InMux I__6015 (
            .O(N__27962),
            .I(N__27914));
    InMux I__6014 (
            .O(N__27959),
            .I(N__27911));
    InMux I__6013 (
            .O(N__27956),
            .I(N__27908));
    LocalMux I__6012 (
            .O(N__27953),
            .I(N__27905));
    LocalMux I__6011 (
            .O(N__27950),
            .I(N__27898));
    Span4Mux_v I__6010 (
            .O(N__27947),
            .I(N__27898));
    LocalMux I__6009 (
            .O(N__27944),
            .I(N__27898));
    LocalMux I__6008 (
            .O(N__27941),
            .I(N__27893));
    Span4Mux_v I__6007 (
            .O(N__27938),
            .I(N__27893));
    Span4Mux_h I__6006 (
            .O(N__27935),
            .I(N__27890));
    Span4Mux_h I__6005 (
            .O(N__27932),
            .I(N__27885));
    Span4Mux_h I__6004 (
            .O(N__27929),
            .I(N__27885));
    Span4Mux_v I__6003 (
            .O(N__27926),
            .I(N__27882));
    Span4Mux_v I__6002 (
            .O(N__27923),
            .I(N__27879));
    Span4Mux_h I__6001 (
            .O(N__27920),
            .I(N__27874));
    Span4Mux_v I__6000 (
            .O(N__27917),
            .I(N__27874));
    LocalMux I__5999 (
            .O(N__27914),
            .I(N__27871));
    LocalMux I__5998 (
            .O(N__27911),
            .I(N__27868));
    LocalMux I__5997 (
            .O(N__27908),
            .I(N__27865));
    Span4Mux_h I__5996 (
            .O(N__27905),
            .I(N__27860));
    Span4Mux_v I__5995 (
            .O(N__27898),
            .I(N__27860));
    Span4Mux_h I__5994 (
            .O(N__27893),
            .I(N__27854));
    Span4Mux_v I__5993 (
            .O(N__27890),
            .I(N__27854));
    Sp12to4 I__5992 (
            .O(N__27885),
            .I(N__27851));
    Sp12to4 I__5991 (
            .O(N__27882),
            .I(N__27844));
    Sp12to4 I__5990 (
            .O(N__27879),
            .I(N__27844));
    Sp12to4 I__5989 (
            .O(N__27874),
            .I(N__27844));
    Span12Mux_h I__5988 (
            .O(N__27871),
            .I(N__27839));
    Span12Mux_h I__5987 (
            .O(N__27868),
            .I(N__27839));
    Span12Mux_h I__5986 (
            .O(N__27865),
            .I(N__27836));
    Span4Mux_h I__5985 (
            .O(N__27860),
            .I(N__27833));
    InMux I__5984 (
            .O(N__27859),
            .I(N__27830));
    Span4Mux_h I__5983 (
            .O(N__27854),
            .I(N__27827));
    Span12Mux_s11_v I__5982 (
            .O(N__27851),
            .I(N__27822));
    Span12Mux_v I__5981 (
            .O(N__27844),
            .I(N__27822));
    Odrv12 I__5980 (
            .O(N__27839),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv12 I__5979 (
            .O(N__27836),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv4 I__5978 (
            .O(N__27833),
            .I(M_this_spr_address_qZ0Z_2));
    LocalMux I__5977 (
            .O(N__27830),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv4 I__5976 (
            .O(N__27827),
            .I(M_this_spr_address_qZ0Z_2));
    Odrv12 I__5975 (
            .O(N__27822),
            .I(M_this_spr_address_qZ0Z_2));
    InMux I__5974 (
            .O(N__27809),
            .I(un1_M_this_spr_address_q_cry_1));
    CascadeMux I__5973 (
            .O(N__27806),
            .I(N__27803));
    InMux I__5972 (
            .O(N__27803),
            .I(N__27799));
    CascadeMux I__5971 (
            .O(N__27802),
            .I(N__27796));
    LocalMux I__5970 (
            .O(N__27799),
            .I(N__27792));
    InMux I__5969 (
            .O(N__27796),
            .I(N__27789));
    CascadeMux I__5968 (
            .O(N__27795),
            .I(N__27786));
    Span4Mux_v I__5967 (
            .O(N__27792),
            .I(N__27779));
    LocalMux I__5966 (
            .O(N__27789),
            .I(N__27779));
    InMux I__5965 (
            .O(N__27786),
            .I(N__27776));
    CascadeMux I__5964 (
            .O(N__27785),
            .I(N__27767));
    CascadeMux I__5963 (
            .O(N__27784),
            .I(N__27764));
    Span4Mux_h I__5962 (
            .O(N__27779),
            .I(N__27757));
    LocalMux I__5961 (
            .O(N__27776),
            .I(N__27757));
    CascadeMux I__5960 (
            .O(N__27775),
            .I(N__27754));
    CascadeMux I__5959 (
            .O(N__27774),
            .I(N__27751));
    CascadeMux I__5958 (
            .O(N__27773),
            .I(N__27748));
    CascadeMux I__5957 (
            .O(N__27772),
            .I(N__27745));
    CascadeMux I__5956 (
            .O(N__27771),
            .I(N__27739));
    CascadeMux I__5955 (
            .O(N__27770),
            .I(N__27736));
    InMux I__5954 (
            .O(N__27767),
            .I(N__27733));
    InMux I__5953 (
            .O(N__27764),
            .I(N__27730));
    CascadeMux I__5952 (
            .O(N__27763),
            .I(N__27727));
    CascadeMux I__5951 (
            .O(N__27762),
            .I(N__27724));
    Span4Mux_v I__5950 (
            .O(N__27757),
            .I(N__27721));
    InMux I__5949 (
            .O(N__27754),
            .I(N__27718));
    InMux I__5948 (
            .O(N__27751),
            .I(N__27715));
    InMux I__5947 (
            .O(N__27748),
            .I(N__27712));
    InMux I__5946 (
            .O(N__27745),
            .I(N__27709));
    CascadeMux I__5945 (
            .O(N__27744),
            .I(N__27706));
    CascadeMux I__5944 (
            .O(N__27743),
            .I(N__27703));
    CascadeMux I__5943 (
            .O(N__27742),
            .I(N__27700));
    InMux I__5942 (
            .O(N__27739),
            .I(N__27697));
    InMux I__5941 (
            .O(N__27736),
            .I(N__27694));
    LocalMux I__5940 (
            .O(N__27733),
            .I(N__27689));
    LocalMux I__5939 (
            .O(N__27730),
            .I(N__27689));
    InMux I__5938 (
            .O(N__27727),
            .I(N__27686));
    InMux I__5937 (
            .O(N__27724),
            .I(N__27683));
    Span4Mux_s1_v I__5936 (
            .O(N__27721),
            .I(N__27678));
    LocalMux I__5935 (
            .O(N__27718),
            .I(N__27678));
    LocalMux I__5934 (
            .O(N__27715),
            .I(N__27675));
    LocalMux I__5933 (
            .O(N__27712),
            .I(N__27672));
    LocalMux I__5932 (
            .O(N__27709),
            .I(N__27669));
    InMux I__5931 (
            .O(N__27706),
            .I(N__27666));
    InMux I__5930 (
            .O(N__27703),
            .I(N__27663));
    InMux I__5929 (
            .O(N__27700),
            .I(N__27660));
    LocalMux I__5928 (
            .O(N__27697),
            .I(N__27657));
    LocalMux I__5927 (
            .O(N__27694),
            .I(N__27652));
    Span4Mux_v I__5926 (
            .O(N__27689),
            .I(N__27652));
    LocalMux I__5925 (
            .O(N__27686),
            .I(N__27647));
    LocalMux I__5924 (
            .O(N__27683),
            .I(N__27647));
    Span4Mux_h I__5923 (
            .O(N__27678),
            .I(N__27644));
    Span4Mux_h I__5922 (
            .O(N__27675),
            .I(N__27641));
    Span4Mux_h I__5921 (
            .O(N__27672),
            .I(N__27638));
    Span4Mux_h I__5920 (
            .O(N__27669),
            .I(N__27635));
    LocalMux I__5919 (
            .O(N__27666),
            .I(N__27632));
    LocalMux I__5918 (
            .O(N__27663),
            .I(N__27629));
    LocalMux I__5917 (
            .O(N__27660),
            .I(N__27626));
    Span4Mux_v I__5916 (
            .O(N__27657),
            .I(N__27619));
    Span4Mux_v I__5915 (
            .O(N__27652),
            .I(N__27619));
    Span4Mux_v I__5914 (
            .O(N__27647),
            .I(N__27619));
    Sp12to4 I__5913 (
            .O(N__27644),
            .I(N__27616));
    Sp12to4 I__5912 (
            .O(N__27641),
            .I(N__27609));
    Sp12to4 I__5911 (
            .O(N__27638),
            .I(N__27609));
    Sp12to4 I__5910 (
            .O(N__27635),
            .I(N__27609));
    Span4Mux_v I__5909 (
            .O(N__27632),
            .I(N__27606));
    Span4Mux_v I__5908 (
            .O(N__27629),
            .I(N__27601));
    Span4Mux_s2_v I__5907 (
            .O(N__27626),
            .I(N__27601));
    Span4Mux_h I__5906 (
            .O(N__27619),
            .I(N__27597));
    Span12Mux_v I__5905 (
            .O(N__27616),
            .I(N__27592));
    Span12Mux_v I__5904 (
            .O(N__27609),
            .I(N__27592));
    Sp12to4 I__5903 (
            .O(N__27606),
            .I(N__27587));
    Sp12to4 I__5902 (
            .O(N__27601),
            .I(N__27587));
    InMux I__5901 (
            .O(N__27600),
            .I(N__27584));
    Span4Mux_h I__5900 (
            .O(N__27597),
            .I(N__27581));
    Span12Mux_h I__5899 (
            .O(N__27592),
            .I(N__27576));
    Span12Mux_h I__5898 (
            .O(N__27587),
            .I(N__27576));
    LocalMux I__5897 (
            .O(N__27584),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv4 I__5896 (
            .O(N__27581),
            .I(M_this_spr_address_qZ0Z_3));
    Odrv12 I__5895 (
            .O(N__27576),
            .I(M_this_spr_address_qZ0Z_3));
    InMux I__5894 (
            .O(N__27569),
            .I(un1_M_this_spr_address_q_cry_2));
    CascadeMux I__5893 (
            .O(N__27566),
            .I(N__27563));
    InMux I__5892 (
            .O(N__27563),
            .I(N__27559));
    CascadeMux I__5891 (
            .O(N__27562),
            .I(N__27556));
    LocalMux I__5890 (
            .O(N__27559),
            .I(N__27547));
    InMux I__5889 (
            .O(N__27556),
            .I(N__27544));
    CascadeMux I__5888 (
            .O(N__27555),
            .I(N__27541));
    CascadeMux I__5887 (
            .O(N__27554),
            .I(N__27537));
    CascadeMux I__5886 (
            .O(N__27553),
            .I(N__27534));
    CascadeMux I__5885 (
            .O(N__27552),
            .I(N__27529));
    CascadeMux I__5884 (
            .O(N__27551),
            .I(N__27526));
    CascadeMux I__5883 (
            .O(N__27550),
            .I(N__27522));
    Span4Mux_s3_v I__5882 (
            .O(N__27547),
            .I(N__27516));
    LocalMux I__5881 (
            .O(N__27544),
            .I(N__27516));
    InMux I__5880 (
            .O(N__27541),
            .I(N__27513));
    CascadeMux I__5879 (
            .O(N__27540),
            .I(N__27510));
    InMux I__5878 (
            .O(N__27537),
            .I(N__27507));
    InMux I__5877 (
            .O(N__27534),
            .I(N__27504));
    CascadeMux I__5876 (
            .O(N__27533),
            .I(N__27501));
    CascadeMux I__5875 (
            .O(N__27532),
            .I(N__27498));
    InMux I__5874 (
            .O(N__27529),
            .I(N__27493));
    InMux I__5873 (
            .O(N__27526),
            .I(N__27490));
    CascadeMux I__5872 (
            .O(N__27525),
            .I(N__27487));
    InMux I__5871 (
            .O(N__27522),
            .I(N__27484));
    CascadeMux I__5870 (
            .O(N__27521),
            .I(N__27481));
    Span4Mux_v I__5869 (
            .O(N__27516),
            .I(N__27476));
    LocalMux I__5868 (
            .O(N__27513),
            .I(N__27476));
    InMux I__5867 (
            .O(N__27510),
            .I(N__27473));
    LocalMux I__5866 (
            .O(N__27507),
            .I(N__27470));
    LocalMux I__5865 (
            .O(N__27504),
            .I(N__27467));
    InMux I__5864 (
            .O(N__27501),
            .I(N__27464));
    InMux I__5863 (
            .O(N__27498),
            .I(N__27460));
    CascadeMux I__5862 (
            .O(N__27497),
            .I(N__27457));
    CascadeMux I__5861 (
            .O(N__27496),
            .I(N__27454));
    LocalMux I__5860 (
            .O(N__27493),
            .I(N__27451));
    LocalMux I__5859 (
            .O(N__27490),
            .I(N__27448));
    InMux I__5858 (
            .O(N__27487),
            .I(N__27445));
    LocalMux I__5857 (
            .O(N__27484),
            .I(N__27442));
    InMux I__5856 (
            .O(N__27481),
            .I(N__27439));
    Span4Mux_h I__5855 (
            .O(N__27476),
            .I(N__27434));
    LocalMux I__5854 (
            .O(N__27473),
            .I(N__27434));
    Span4Mux_v I__5853 (
            .O(N__27470),
            .I(N__27427));
    Span4Mux_h I__5852 (
            .O(N__27467),
            .I(N__27427));
    LocalMux I__5851 (
            .O(N__27464),
            .I(N__27427));
    CascadeMux I__5850 (
            .O(N__27463),
            .I(N__27424));
    LocalMux I__5849 (
            .O(N__27460),
            .I(N__27421));
    InMux I__5848 (
            .O(N__27457),
            .I(N__27418));
    InMux I__5847 (
            .O(N__27454),
            .I(N__27415));
    Span4Mux_v I__5846 (
            .O(N__27451),
            .I(N__27410));
    Span4Mux_h I__5845 (
            .O(N__27448),
            .I(N__27410));
    LocalMux I__5844 (
            .O(N__27445),
            .I(N__27407));
    Span4Mux_h I__5843 (
            .O(N__27442),
            .I(N__27402));
    LocalMux I__5842 (
            .O(N__27439),
            .I(N__27402));
    Span4Mux_v I__5841 (
            .O(N__27434),
            .I(N__27397));
    Span4Mux_v I__5840 (
            .O(N__27427),
            .I(N__27397));
    InMux I__5839 (
            .O(N__27424),
            .I(N__27394));
    Span12Mux_h I__5838 (
            .O(N__27421),
            .I(N__27391));
    LocalMux I__5837 (
            .O(N__27418),
            .I(N__27388));
    LocalMux I__5836 (
            .O(N__27415),
            .I(N__27385));
    Sp12to4 I__5835 (
            .O(N__27410),
            .I(N__27382));
    Sp12to4 I__5834 (
            .O(N__27407),
            .I(N__27377));
    Sp12to4 I__5833 (
            .O(N__27402),
            .I(N__27377));
    Sp12to4 I__5832 (
            .O(N__27397),
            .I(N__27372));
    LocalMux I__5831 (
            .O(N__27394),
            .I(N__27372));
    Span12Mux_v I__5830 (
            .O(N__27391),
            .I(N__27364));
    Span12Mux_h I__5829 (
            .O(N__27388),
            .I(N__27364));
    Span12Mux_h I__5828 (
            .O(N__27385),
            .I(N__27364));
    Span12Mux_v I__5827 (
            .O(N__27382),
            .I(N__27357));
    Span12Mux_s11_v I__5826 (
            .O(N__27377),
            .I(N__27357));
    Span12Mux_s11_h I__5825 (
            .O(N__27372),
            .I(N__27357));
    InMux I__5824 (
            .O(N__27371),
            .I(N__27354));
    Odrv12 I__5823 (
            .O(N__27364),
            .I(M_this_spr_address_qZ0Z_4));
    Odrv12 I__5822 (
            .O(N__27357),
            .I(M_this_spr_address_qZ0Z_4));
    LocalMux I__5821 (
            .O(N__27354),
            .I(M_this_spr_address_qZ0Z_4));
    InMux I__5820 (
            .O(N__27347),
            .I(un1_M_this_spr_address_q_cry_3));
    CascadeMux I__5819 (
            .O(N__27344),
            .I(N__27340));
    CascadeMux I__5818 (
            .O(N__27343),
            .I(N__27337));
    InMux I__5817 (
            .O(N__27340),
            .I(N__27330));
    InMux I__5816 (
            .O(N__27337),
            .I(N__27327));
    CascadeMux I__5815 (
            .O(N__27336),
            .I(N__27324));
    CascadeMux I__5814 (
            .O(N__27335),
            .I(N__27321));
    CascadeMux I__5813 (
            .O(N__27334),
            .I(N__27313));
    CascadeMux I__5812 (
            .O(N__27333),
            .I(N__27309));
    LocalMux I__5811 (
            .O(N__27330),
            .I(N__27304));
    LocalMux I__5810 (
            .O(N__27327),
            .I(N__27304));
    InMux I__5809 (
            .O(N__27324),
            .I(N__27301));
    InMux I__5808 (
            .O(N__27321),
            .I(N__27298));
    CascadeMux I__5807 (
            .O(N__27320),
            .I(N__27295));
    CascadeMux I__5806 (
            .O(N__27319),
            .I(N__27292));
    CascadeMux I__5805 (
            .O(N__27318),
            .I(N__27289));
    CascadeMux I__5804 (
            .O(N__27317),
            .I(N__27286));
    CascadeMux I__5803 (
            .O(N__27316),
            .I(N__27283));
    InMux I__5802 (
            .O(N__27313),
            .I(N__27277));
    CascadeMux I__5801 (
            .O(N__27312),
            .I(N__27273));
    InMux I__5800 (
            .O(N__27309),
            .I(N__27270));
    Span4Mux_v I__5799 (
            .O(N__27304),
            .I(N__27263));
    LocalMux I__5798 (
            .O(N__27301),
            .I(N__27263));
    LocalMux I__5797 (
            .O(N__27298),
            .I(N__27263));
    InMux I__5796 (
            .O(N__27295),
            .I(N__27260));
    InMux I__5795 (
            .O(N__27292),
            .I(N__27257));
    InMux I__5794 (
            .O(N__27289),
            .I(N__27254));
    InMux I__5793 (
            .O(N__27286),
            .I(N__27251));
    InMux I__5792 (
            .O(N__27283),
            .I(N__27248));
    CascadeMux I__5791 (
            .O(N__27282),
            .I(N__27245));
    CascadeMux I__5790 (
            .O(N__27281),
            .I(N__27242));
    CascadeMux I__5789 (
            .O(N__27280),
            .I(N__27239));
    LocalMux I__5788 (
            .O(N__27277),
            .I(N__27236));
    CascadeMux I__5787 (
            .O(N__27276),
            .I(N__27233));
    InMux I__5786 (
            .O(N__27273),
            .I(N__27230));
    LocalMux I__5785 (
            .O(N__27270),
            .I(N__27227));
    Span4Mux_v I__5784 (
            .O(N__27263),
            .I(N__27222));
    LocalMux I__5783 (
            .O(N__27260),
            .I(N__27222));
    LocalMux I__5782 (
            .O(N__27257),
            .I(N__27217));
    LocalMux I__5781 (
            .O(N__27254),
            .I(N__27217));
    LocalMux I__5780 (
            .O(N__27251),
            .I(N__27212));
    LocalMux I__5779 (
            .O(N__27248),
            .I(N__27212));
    InMux I__5778 (
            .O(N__27245),
            .I(N__27209));
    InMux I__5777 (
            .O(N__27242),
            .I(N__27206));
    InMux I__5776 (
            .O(N__27239),
            .I(N__27203));
    Span4Mux_v I__5775 (
            .O(N__27236),
            .I(N__27200));
    InMux I__5774 (
            .O(N__27233),
            .I(N__27197));
    LocalMux I__5773 (
            .O(N__27230),
            .I(N__27194));
    Span4Mux_v I__5772 (
            .O(N__27227),
            .I(N__27191));
    Span4Mux_v I__5771 (
            .O(N__27222),
            .I(N__27188));
    Span4Mux_v I__5770 (
            .O(N__27217),
            .I(N__27183));
    Span4Mux_v I__5769 (
            .O(N__27212),
            .I(N__27183));
    LocalMux I__5768 (
            .O(N__27209),
            .I(N__27175));
    LocalMux I__5767 (
            .O(N__27206),
            .I(N__27175));
    LocalMux I__5766 (
            .O(N__27203),
            .I(N__27175));
    Sp12to4 I__5765 (
            .O(N__27200),
            .I(N__27166));
    LocalMux I__5764 (
            .O(N__27197),
            .I(N__27166));
    Span12Mux_s8_v I__5763 (
            .O(N__27194),
            .I(N__27166));
    Sp12to4 I__5762 (
            .O(N__27191),
            .I(N__27166));
    Sp12to4 I__5761 (
            .O(N__27188),
            .I(N__27163));
    Sp12to4 I__5760 (
            .O(N__27183),
            .I(N__27160));
    InMux I__5759 (
            .O(N__27182),
            .I(N__27157));
    Span12Mux_s11_v I__5758 (
            .O(N__27175),
            .I(N__27152));
    Span12Mux_v I__5757 (
            .O(N__27166),
            .I(N__27152));
    Span12Mux_h I__5756 (
            .O(N__27163),
            .I(N__27147));
    Span12Mux_h I__5755 (
            .O(N__27160),
            .I(N__27147));
    LocalMux I__5754 (
            .O(N__27157),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv12 I__5753 (
            .O(N__27152),
            .I(M_this_spr_address_qZ0Z_5));
    Odrv12 I__5752 (
            .O(N__27147),
            .I(M_this_spr_address_qZ0Z_5));
    InMux I__5751 (
            .O(N__27140),
            .I(un1_M_this_spr_address_q_cry_4));
    CascadeMux I__5750 (
            .O(N__27137),
            .I(N__27131));
    CascadeMux I__5749 (
            .O(N__27136),
            .I(N__27127));
    CascadeMux I__5748 (
            .O(N__27135),
            .I(N__27124));
    CascadeMux I__5747 (
            .O(N__27134),
            .I(N__27121));
    InMux I__5746 (
            .O(N__27131),
            .I(N__27117));
    CascadeMux I__5745 (
            .O(N__27130),
            .I(N__27114));
    InMux I__5744 (
            .O(N__27127),
            .I(N__27110));
    InMux I__5743 (
            .O(N__27124),
            .I(N__27107));
    InMux I__5742 (
            .O(N__27121),
            .I(N__27102));
    CascadeMux I__5741 (
            .O(N__27120),
            .I(N__27099));
    LocalMux I__5740 (
            .O(N__27117),
            .I(N__27096));
    InMux I__5739 (
            .O(N__27114),
            .I(N__27093));
    CascadeMux I__5738 (
            .O(N__27113),
            .I(N__27090));
    LocalMux I__5737 (
            .O(N__27110),
            .I(N__27087));
    LocalMux I__5736 (
            .O(N__27107),
            .I(N__27084));
    CascadeMux I__5735 (
            .O(N__27106),
            .I(N__27080));
    CascadeMux I__5734 (
            .O(N__27105),
            .I(N__27076));
    LocalMux I__5733 (
            .O(N__27102),
            .I(N__27070));
    InMux I__5732 (
            .O(N__27099),
            .I(N__27067));
    Span4Mux_s2_v I__5731 (
            .O(N__27096),
            .I(N__27061));
    LocalMux I__5730 (
            .O(N__27093),
            .I(N__27061));
    InMux I__5729 (
            .O(N__27090),
            .I(N__27058));
    Span4Mux_h I__5728 (
            .O(N__27087),
            .I(N__27055));
    Span4Mux_h I__5727 (
            .O(N__27084),
            .I(N__27052));
    CascadeMux I__5726 (
            .O(N__27083),
            .I(N__27049));
    InMux I__5725 (
            .O(N__27080),
            .I(N__27046));
    CascadeMux I__5724 (
            .O(N__27079),
            .I(N__27043));
    InMux I__5723 (
            .O(N__27076),
            .I(N__27040));
    CascadeMux I__5722 (
            .O(N__27075),
            .I(N__27037));
    CascadeMux I__5721 (
            .O(N__27074),
            .I(N__27034));
    CascadeMux I__5720 (
            .O(N__27073),
            .I(N__27030));
    Span4Mux_h I__5719 (
            .O(N__27070),
            .I(N__27025));
    LocalMux I__5718 (
            .O(N__27067),
            .I(N__27025));
    CascadeMux I__5717 (
            .O(N__27066),
            .I(N__27022));
    Span4Mux_v I__5716 (
            .O(N__27061),
            .I(N__27017));
    LocalMux I__5715 (
            .O(N__27058),
            .I(N__27017));
    Span4Mux_h I__5714 (
            .O(N__27055),
            .I(N__27014));
    Span4Mux_h I__5713 (
            .O(N__27052),
            .I(N__27011));
    InMux I__5712 (
            .O(N__27049),
            .I(N__27008));
    LocalMux I__5711 (
            .O(N__27046),
            .I(N__27005));
    InMux I__5710 (
            .O(N__27043),
            .I(N__27002));
    LocalMux I__5709 (
            .O(N__27040),
            .I(N__26999));
    InMux I__5708 (
            .O(N__27037),
            .I(N__26996));
    InMux I__5707 (
            .O(N__27034),
            .I(N__26993));
    CascadeMux I__5706 (
            .O(N__27033),
            .I(N__26990));
    InMux I__5705 (
            .O(N__27030),
            .I(N__26987));
    Span4Mux_v I__5704 (
            .O(N__27025),
            .I(N__26984));
    InMux I__5703 (
            .O(N__27022),
            .I(N__26981));
    Span4Mux_v I__5702 (
            .O(N__27017),
            .I(N__26978));
    Span4Mux_v I__5701 (
            .O(N__27014),
            .I(N__26975));
    Span4Mux_v I__5700 (
            .O(N__27011),
            .I(N__26972));
    LocalMux I__5699 (
            .O(N__27008),
            .I(N__26969));
    Span4Mux_h I__5698 (
            .O(N__27005),
            .I(N__26964));
    LocalMux I__5697 (
            .O(N__27002),
            .I(N__26964));
    Span4Mux_v I__5696 (
            .O(N__26999),
            .I(N__26957));
    LocalMux I__5695 (
            .O(N__26996),
            .I(N__26957));
    LocalMux I__5694 (
            .O(N__26993),
            .I(N__26957));
    InMux I__5693 (
            .O(N__26990),
            .I(N__26954));
    LocalMux I__5692 (
            .O(N__26987),
            .I(N__26951));
    Sp12to4 I__5691 (
            .O(N__26984),
            .I(N__26946));
    LocalMux I__5690 (
            .O(N__26981),
            .I(N__26946));
    Span4Mux_h I__5689 (
            .O(N__26978),
            .I(N__26943));
    Sp12to4 I__5688 (
            .O(N__26975),
            .I(N__26936));
    Sp12to4 I__5687 (
            .O(N__26972),
            .I(N__26936));
    Span12Mux_h I__5686 (
            .O(N__26969),
            .I(N__26936));
    Span4Mux_v I__5685 (
            .O(N__26964),
            .I(N__26929));
    Span4Mux_v I__5684 (
            .O(N__26957),
            .I(N__26929));
    LocalMux I__5683 (
            .O(N__26954),
            .I(N__26929));
    Span12Mux_h I__5682 (
            .O(N__26951),
            .I(N__26923));
    Span12Mux_h I__5681 (
            .O(N__26946),
            .I(N__26923));
    Span4Mux_h I__5680 (
            .O(N__26943),
            .I(N__26920));
    Span12Mux_v I__5679 (
            .O(N__26936),
            .I(N__26915));
    Sp12to4 I__5678 (
            .O(N__26929),
            .I(N__26915));
    InMux I__5677 (
            .O(N__26928),
            .I(N__26912));
    Odrv12 I__5676 (
            .O(N__26923),
            .I(M_this_spr_address_qZ0Z_6));
    Odrv4 I__5675 (
            .O(N__26920),
            .I(M_this_spr_address_qZ0Z_6));
    Odrv12 I__5674 (
            .O(N__26915),
            .I(M_this_spr_address_qZ0Z_6));
    LocalMux I__5673 (
            .O(N__26912),
            .I(M_this_spr_address_qZ0Z_6));
    InMux I__5672 (
            .O(N__26903),
            .I(un1_M_this_spr_address_q_cry_5));
    InMux I__5671 (
            .O(N__26900),
            .I(N__26897));
    LocalMux I__5670 (
            .O(N__26897),
            .I(M_this_data_count_q_cry_11_THRU_CO));
    InMux I__5669 (
            .O(N__26894),
            .I(N__26891));
    LocalMux I__5668 (
            .O(N__26891),
            .I(M_this_data_count_q_s_13));
    InMux I__5667 (
            .O(N__26888),
            .I(N__26885));
    LocalMux I__5666 (
            .O(N__26885),
            .I(M_this_data_count_q_cry_10_THRU_CO));
    InMux I__5665 (
            .O(N__26882),
            .I(N__26877));
    InMux I__5664 (
            .O(N__26881),
            .I(N__26874));
    InMux I__5663 (
            .O(N__26880),
            .I(N__26871));
    LocalMux I__5662 (
            .O(N__26877),
            .I(N__26868));
    LocalMux I__5661 (
            .O(N__26874),
            .I(N__26865));
    LocalMux I__5660 (
            .O(N__26871),
            .I(M_this_data_count_qZ0Z_7));
    Odrv4 I__5659 (
            .O(N__26868),
            .I(M_this_data_count_qZ0Z_7));
    Odrv4 I__5658 (
            .O(N__26865),
            .I(M_this_data_count_qZ0Z_7));
    InMux I__5657 (
            .O(N__26858),
            .I(N__26855));
    LocalMux I__5656 (
            .O(N__26855),
            .I(N__26852));
    Odrv4 I__5655 (
            .O(N__26852),
            .I(\this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11 ));
    CascadeMux I__5654 (
            .O(N__26849),
            .I(\this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_ ));
    InMux I__5653 (
            .O(N__26846),
            .I(N__26843));
    LocalMux I__5652 (
            .O(N__26843),
            .I(\this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11 ));
    InMux I__5651 (
            .O(N__26840),
            .I(N__26835));
    InMux I__5650 (
            .O(N__26839),
            .I(N__26830));
    InMux I__5649 (
            .O(N__26838),
            .I(N__26830));
    LocalMux I__5648 (
            .O(N__26835),
            .I(M_this_data_count_qZ0Z_12));
    LocalMux I__5647 (
            .O(N__26830),
            .I(M_this_data_count_qZ0Z_12));
    CascadeMux I__5646 (
            .O(N__26825),
            .I(N__26822));
    InMux I__5645 (
            .O(N__26822),
            .I(N__26817));
    InMux I__5644 (
            .O(N__26821),
            .I(N__26812));
    InMux I__5643 (
            .O(N__26820),
            .I(N__26812));
    LocalMux I__5642 (
            .O(N__26817),
            .I(M_this_data_count_qZ0Z_11));
    LocalMux I__5641 (
            .O(N__26812),
            .I(M_this_data_count_qZ0Z_11));
    CascadeMux I__5640 (
            .O(N__26807),
            .I(N__26803));
    InMux I__5639 (
            .O(N__26806),
            .I(N__26800));
    InMux I__5638 (
            .O(N__26803),
            .I(N__26797));
    LocalMux I__5637 (
            .O(N__26800),
            .I(M_this_data_count_qZ0Z_13));
    LocalMux I__5636 (
            .O(N__26797),
            .I(M_this_data_count_qZ0Z_13));
    InMux I__5635 (
            .O(N__26792),
            .I(N__26788));
    InMux I__5634 (
            .O(N__26791),
            .I(N__26785));
    LocalMux I__5633 (
            .O(N__26788),
            .I(M_this_data_count_qZ0Z_10));
    LocalMux I__5632 (
            .O(N__26785),
            .I(M_this_data_count_qZ0Z_10));
    InMux I__5631 (
            .O(N__26780),
            .I(N__26777));
    LocalMux I__5630 (
            .O(N__26777),
            .I(\this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11 ));
    CascadeMux I__5629 (
            .O(N__26774),
            .I(N__26771));
    InMux I__5628 (
            .O(N__26771),
            .I(N__26768));
    LocalMux I__5627 (
            .O(N__26768),
            .I(N__26765));
    Odrv4 I__5626 (
            .O(N__26765),
            .I(M_this_data_count_q_cry_5_THRU_CO));
    InMux I__5625 (
            .O(N__26762),
            .I(N__26741));
    InMux I__5624 (
            .O(N__26761),
            .I(N__26741));
    InMux I__5623 (
            .O(N__26760),
            .I(N__26741));
    InMux I__5622 (
            .O(N__26759),
            .I(N__26741));
    InMux I__5621 (
            .O(N__26758),
            .I(N__26730));
    InMux I__5620 (
            .O(N__26757),
            .I(N__26730));
    InMux I__5619 (
            .O(N__26756),
            .I(N__26730));
    InMux I__5618 (
            .O(N__26755),
            .I(N__26730));
    InMux I__5617 (
            .O(N__26754),
            .I(N__26730));
    InMux I__5616 (
            .O(N__26753),
            .I(N__26721));
    InMux I__5615 (
            .O(N__26752),
            .I(N__26721));
    InMux I__5614 (
            .O(N__26751),
            .I(N__26721));
    InMux I__5613 (
            .O(N__26750),
            .I(N__26721));
    LocalMux I__5612 (
            .O(N__26741),
            .I(N_685_i));
    LocalMux I__5611 (
            .O(N__26730),
            .I(N_685_i));
    LocalMux I__5610 (
            .O(N__26721),
            .I(N_685_i));
    CascadeMux I__5609 (
            .O(N__26714),
            .I(N__26711));
    InMux I__5608 (
            .O(N__26711),
            .I(N__26708));
    LocalMux I__5607 (
            .O(N__26708),
            .I(N__26705));
    Sp12to4 I__5606 (
            .O(N__26705),
            .I(N__26700));
    InMux I__5605 (
            .O(N__26704),
            .I(N__26695));
    InMux I__5604 (
            .O(N__26703),
            .I(N__26695));
    Odrv12 I__5603 (
            .O(N__26700),
            .I(M_this_data_count_qZ0Z_6));
    LocalMux I__5602 (
            .O(N__26695),
            .I(M_this_data_count_qZ0Z_6));
    InMux I__5601 (
            .O(N__26690),
            .I(N__26687));
    LocalMux I__5600 (
            .O(N__26687),
            .I(N__26684));
    Span4Mux_h I__5599 (
            .O(N__26684),
            .I(N__26680));
    InMux I__5598 (
            .O(N__26683),
            .I(N__26677));
    Span4Mux_v I__5597 (
            .O(N__26680),
            .I(N__26674));
    LocalMux I__5596 (
            .O(N__26677),
            .I(M_this_ctrl_flags_qZ0Z_5));
    Odrv4 I__5595 (
            .O(N__26674),
            .I(M_this_ctrl_flags_qZ0Z_5));
    InMux I__5594 (
            .O(N__26669),
            .I(N__26663));
    InMux I__5593 (
            .O(N__26668),
            .I(N__26660));
    InMux I__5592 (
            .O(N__26667),
            .I(N__26656));
    InMux I__5591 (
            .O(N__26666),
            .I(N__26653));
    LocalMux I__5590 (
            .O(N__26663),
            .I(N__26648));
    LocalMux I__5589 (
            .O(N__26660),
            .I(N__26648));
    InMux I__5588 (
            .O(N__26659),
            .I(N__26645));
    LocalMux I__5587 (
            .O(N__26656),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__5586 (
            .O(N__26653),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    Odrv12 I__5585 (
            .O(N__26648),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    LocalMux I__5584 (
            .O(N__26645),
            .I(\this_vga_signals.M_vcounter_qZ0Z_1 ));
    CascadeMux I__5583 (
            .O(N__26636),
            .I(\this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_ ));
    InMux I__5582 (
            .O(N__26633),
            .I(N__26630));
    LocalMux I__5581 (
            .O(N__26630),
            .I(\this_vga_signals.g0_i_x2_4 ));
    CascadeMux I__5580 (
            .O(N__26627),
            .I(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_ ));
    CascadeMux I__5579 (
            .O(N__26624),
            .I(N__26621));
    InMux I__5578 (
            .O(N__26621),
            .I(N__26618));
    LocalMux I__5577 (
            .O(N__26618),
            .I(\this_vga_signals.N_17_i ));
    InMux I__5576 (
            .O(N__26615),
            .I(N__26612));
    LocalMux I__5575 (
            .O(N__26612),
            .I(M_this_data_count_q_s_10));
    InMux I__5574 (
            .O(N__26609),
            .I(N__26606));
    LocalMux I__5573 (
            .O(N__26606),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_11 ));
    InMux I__5572 (
            .O(N__26603),
            .I(N__26600));
    LocalMux I__5571 (
            .O(N__26600),
            .I(N__26597));
    Span12Mux_h I__5570 (
            .O(N__26597),
            .I(N__26594));
    Odrv12 I__5569 (
            .O(N__26594),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_12 ));
    InMux I__5568 (
            .O(N__26591),
            .I(N__26588));
    LocalMux I__5567 (
            .O(N__26588),
            .I(\this_ppu.M_oam_cache_read_data_i_12 ));
    InMux I__5566 (
            .O(N__26585),
            .I(N__26582));
    LocalMux I__5565 (
            .O(N__26582),
            .I(N__26579));
    Span4Mux_h I__5564 (
            .O(N__26579),
            .I(N__26576));
    Span4Mux_h I__5563 (
            .O(N__26576),
            .I(N__26573));
    Span4Mux_h I__5562 (
            .O(N__26573),
            .I(N__26570));
    Odrv4 I__5561 (
            .O(N__26570),
            .I(\this_ppu.oam_cache.mem_8 ));
    CascadeMux I__5560 (
            .O(N__26567),
            .I(N__26564));
    InMux I__5559 (
            .O(N__26564),
            .I(N__26561));
    LocalMux I__5558 (
            .O(N__26561),
            .I(N__26558));
    Span4Mux_v I__5557 (
            .O(N__26558),
            .I(N__26555));
    Span4Mux_h I__5556 (
            .O(N__26555),
            .I(N__26551));
    InMux I__5555 (
            .O(N__26554),
            .I(N__26548));
    Odrv4 I__5554 (
            .O(N__26551),
            .I(\this_ppu.M_oam_cache_read_data_8 ));
    LocalMux I__5553 (
            .O(N__26548),
            .I(\this_ppu.M_oam_cache_read_data_8 ));
    InMux I__5552 (
            .O(N__26543),
            .I(N__26540));
    LocalMux I__5551 (
            .O(N__26540),
            .I(N__26537));
    Span4Mux_v I__5550 (
            .O(N__26537),
            .I(N__26532));
    InMux I__5549 (
            .O(N__26536),
            .I(N__26529));
    InMux I__5548 (
            .O(N__26535),
            .I(N__26526));
    Odrv4 I__5547 (
            .O(N__26532),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__5546 (
            .O(N__26529),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    LocalMux I__5545 (
            .O(N__26526),
            .I(\this_vga_signals.M_vcounter_qZ0Z_0 ));
    CascadeMux I__5544 (
            .O(N__26519),
            .I(\this_vga_signals.N_3_1_cascade_ ));
    InMux I__5543 (
            .O(N__26516),
            .I(N__26513));
    LocalMux I__5542 (
            .O(N__26513),
            .I(N__26510));
    Odrv4 I__5541 (
            .O(N__26510),
            .I(\this_vga_signals.g0_41_N_2L1 ));
    CascadeMux I__5540 (
            .O(N__26507),
            .I(\this_vga_signals.g0_41_N_4L5_cascade_ ));
    InMux I__5539 (
            .O(N__26504),
            .I(N__26501));
    LocalMux I__5538 (
            .O(N__26501),
            .I(\this_vga_signals.g0_41_1 ));
    CascadeMux I__5537 (
            .O(N__26498),
            .I(N__26495));
    InMux I__5536 (
            .O(N__26495),
            .I(N__26492));
    LocalMux I__5535 (
            .O(N__26492),
            .I(N__26488));
    InMux I__5534 (
            .O(N__26491),
            .I(N__26485));
    Span4Mux_v I__5533 (
            .O(N__26488),
            .I(N__26482));
    LocalMux I__5532 (
            .O(N__26485),
            .I(N__26475));
    Span4Mux_h I__5531 (
            .O(N__26482),
            .I(N__26475));
    InMux I__5530 (
            .O(N__26481),
            .I(N__26470));
    InMux I__5529 (
            .O(N__26480),
            .I(N__26470));
    Span4Mux_h I__5528 (
            .O(N__26475),
            .I(N__26463));
    LocalMux I__5527 (
            .O(N__26470),
            .I(N__26463));
    InMux I__5526 (
            .O(N__26469),
            .I(N__26457));
    InMux I__5525 (
            .O(N__26468),
            .I(N__26454));
    Span4Mux_h I__5524 (
            .O(N__26463),
            .I(N__26451));
    InMux I__5523 (
            .O(N__26462),
            .I(N__26444));
    InMux I__5522 (
            .O(N__26461),
            .I(N__26444));
    InMux I__5521 (
            .O(N__26460),
            .I(N__26444));
    LocalMux I__5520 (
            .O(N__26457),
            .I(N__26439));
    LocalMux I__5519 (
            .O(N__26454),
            .I(N__26439));
    Odrv4 I__5518 (
            .O(N__26451),
            .I(M_this_vga_ramdac_en));
    LocalMux I__5517 (
            .O(N__26444),
            .I(M_this_vga_ramdac_en));
    Odrv4 I__5516 (
            .O(N__26439),
            .I(M_this_vga_ramdac_en));
    InMux I__5515 (
            .O(N__26432),
            .I(N__26429));
    LocalMux I__5514 (
            .O(N__26429),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_0_0_1 ));
    CascadeMux I__5513 (
            .O(N__26426),
            .I(N__26423));
    InMux I__5512 (
            .O(N__26423),
            .I(N__26420));
    LocalMux I__5511 (
            .O(N__26420),
            .I(N__26417));
    Span4Mux_h I__5510 (
            .O(N__26417),
            .I(N__26414));
    Span4Mux_h I__5509 (
            .O(N__26414),
            .I(N__26411));
    Odrv4 I__5508 (
            .O(N__26411),
            .I(M_this_vga_signals_address_7));
    InMux I__5507 (
            .O(N__26408),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_4 ));
    InMux I__5506 (
            .O(N__26405),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_5 ));
    InMux I__5505 (
            .O(N__26402),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_6 ));
    InMux I__5504 (
            .O(N__26399),
            .I(bfn_16_16_0_));
    InMux I__5503 (
            .O(N__26396),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_8 ));
    InMux I__5502 (
            .O(N__26393),
            .I(N__26390));
    LocalMux I__5501 (
            .O(N__26390),
            .I(\this_vga_signals.M_vcounter_d7lto9_i_a2_1 ));
    IoInMux I__5500 (
            .O(N__26387),
            .I(N__26384));
    LocalMux I__5499 (
            .O(N__26384),
            .I(N__26381));
    Span4Mux_s3_h I__5498 (
            .O(N__26381),
            .I(N__26378));
    Span4Mux_h I__5497 (
            .O(N__26378),
            .I(N__26375));
    Span4Mux_h I__5496 (
            .O(N__26375),
            .I(N__26372));
    Span4Mux_h I__5495 (
            .O(N__26372),
            .I(N__26369));
    Span4Mux_v I__5494 (
            .O(N__26369),
            .I(N__26366));
    Odrv4 I__5493 (
            .O(N__26366),
            .I(port_nmib_1_i));
    InMux I__5492 (
            .O(N__26363),
            .I(N__26360));
    LocalMux I__5491 (
            .O(N__26360),
            .I(\this_ppu.M_oam_cache_read_data_i_11 ));
    InMux I__5490 (
            .O(N__26357),
            .I(N__26354));
    LocalMux I__5489 (
            .O(N__26354),
            .I(N__26351));
    Span4Mux_h I__5488 (
            .O(N__26351),
            .I(N__26348));
    Span4Mux_h I__5487 (
            .O(N__26348),
            .I(N__26345));
    Odrv4 I__5486 (
            .O(N__26345),
            .I(\this_ppu.oam_cache.mem_11 ));
    InMux I__5485 (
            .O(N__26342),
            .I(N__26339));
    LocalMux I__5484 (
            .O(N__26339),
            .I(\this_reset_cond.M_stage_qZ0Z_3 ));
    InMux I__5483 (
            .O(N__26336),
            .I(N__26333));
    LocalMux I__5482 (
            .O(N__26333),
            .I(\this_reset_cond.M_stage_qZ0Z_4 ));
    InMux I__5481 (
            .O(N__26330),
            .I(N__26327));
    LocalMux I__5480 (
            .O(N__26327),
            .I(\this_reset_cond.M_stage_qZ0Z_0 ));
    InMux I__5479 (
            .O(N__26324),
            .I(N__26321));
    LocalMux I__5478 (
            .O(N__26321),
            .I(N__26318));
    Span4Mux_v I__5477 (
            .O(N__26318),
            .I(N__26315));
    Span4Mux_v I__5476 (
            .O(N__26315),
            .I(N__26312));
    Span4Mux_v I__5475 (
            .O(N__26312),
            .I(N__26309));
    Span4Mux_h I__5474 (
            .O(N__26309),
            .I(N__26306));
    Span4Mux_h I__5473 (
            .O(N__26306),
            .I(N__26303));
    Odrv4 I__5472 (
            .O(N__26303),
            .I(M_this_map_ram_read_data_0));
    CascadeMux I__5471 (
            .O(N__26300),
            .I(N__26291));
    CascadeMux I__5470 (
            .O(N__26299),
            .I(N__26286));
    CascadeMux I__5469 (
            .O(N__26298),
            .I(N__26283));
    CascadeMux I__5468 (
            .O(N__26297),
            .I(N__26280));
    CascadeMux I__5467 (
            .O(N__26296),
            .I(N__26273));
    CascadeMux I__5466 (
            .O(N__26295),
            .I(N__26270));
    CascadeMux I__5465 (
            .O(N__26294),
            .I(N__26267));
    InMux I__5464 (
            .O(N__26291),
            .I(N__26264));
    CascadeMux I__5463 (
            .O(N__26290),
            .I(N__26260));
    CascadeMux I__5462 (
            .O(N__26289),
            .I(N__26257));
    InMux I__5461 (
            .O(N__26286),
            .I(N__26254));
    InMux I__5460 (
            .O(N__26283),
            .I(N__26251));
    InMux I__5459 (
            .O(N__26280),
            .I(N__26248));
    CascadeMux I__5458 (
            .O(N__26279),
            .I(N__26245));
    CascadeMux I__5457 (
            .O(N__26278),
            .I(N__26242));
    CascadeMux I__5456 (
            .O(N__26277),
            .I(N__26239));
    CascadeMux I__5455 (
            .O(N__26276),
            .I(N__26236));
    InMux I__5454 (
            .O(N__26273),
            .I(N__26233));
    InMux I__5453 (
            .O(N__26270),
            .I(N__26230));
    InMux I__5452 (
            .O(N__26267),
            .I(N__26227));
    LocalMux I__5451 (
            .O(N__26264),
            .I(N__26224));
    CascadeMux I__5450 (
            .O(N__26263),
            .I(N__26221));
    InMux I__5449 (
            .O(N__26260),
            .I(N__26216));
    InMux I__5448 (
            .O(N__26257),
            .I(N__26213));
    LocalMux I__5447 (
            .O(N__26254),
            .I(N__26210));
    LocalMux I__5446 (
            .O(N__26251),
            .I(N__26207));
    LocalMux I__5445 (
            .O(N__26248),
            .I(N__26204));
    InMux I__5444 (
            .O(N__26245),
            .I(N__26201));
    InMux I__5443 (
            .O(N__26242),
            .I(N__26198));
    InMux I__5442 (
            .O(N__26239),
            .I(N__26195));
    InMux I__5441 (
            .O(N__26236),
            .I(N__26192));
    LocalMux I__5440 (
            .O(N__26233),
            .I(N__26189));
    LocalMux I__5439 (
            .O(N__26230),
            .I(N__26186));
    LocalMux I__5438 (
            .O(N__26227),
            .I(N__26183));
    Span4Mux_v I__5437 (
            .O(N__26224),
            .I(N__26180));
    InMux I__5436 (
            .O(N__26221),
            .I(N__26177));
    CascadeMux I__5435 (
            .O(N__26220),
            .I(N__26174));
    CascadeMux I__5434 (
            .O(N__26219),
            .I(N__26171));
    LocalMux I__5433 (
            .O(N__26216),
            .I(N__26168));
    LocalMux I__5432 (
            .O(N__26213),
            .I(N__26165));
    Span4Mux_h I__5431 (
            .O(N__26210),
            .I(N__26162));
    Span4Mux_h I__5430 (
            .O(N__26207),
            .I(N__26159));
    Span4Mux_h I__5429 (
            .O(N__26204),
            .I(N__26156));
    LocalMux I__5428 (
            .O(N__26201),
            .I(N__26153));
    LocalMux I__5427 (
            .O(N__26198),
            .I(N__26148));
    LocalMux I__5426 (
            .O(N__26195),
            .I(N__26148));
    LocalMux I__5425 (
            .O(N__26192),
            .I(N__26141));
    Span4Mux_h I__5424 (
            .O(N__26189),
            .I(N__26141));
    Span4Mux_v I__5423 (
            .O(N__26186),
            .I(N__26141));
    Sp12to4 I__5422 (
            .O(N__26183),
            .I(N__26138));
    Sp12to4 I__5421 (
            .O(N__26180),
            .I(N__26133));
    LocalMux I__5420 (
            .O(N__26177),
            .I(N__26133));
    InMux I__5419 (
            .O(N__26174),
            .I(N__26130));
    InMux I__5418 (
            .O(N__26171),
            .I(N__26127));
    Span4Mux_h I__5417 (
            .O(N__26168),
            .I(N__26124));
    Span4Mux_h I__5416 (
            .O(N__26165),
            .I(N__26121));
    Span4Mux_h I__5415 (
            .O(N__26162),
            .I(N__26118));
    Span4Mux_h I__5414 (
            .O(N__26159),
            .I(N__26113));
    Span4Mux_h I__5413 (
            .O(N__26156),
            .I(N__26113));
    Span4Mux_h I__5412 (
            .O(N__26153),
            .I(N__26106));
    Span4Mux_v I__5411 (
            .O(N__26148),
            .I(N__26106));
    Span4Mux_v I__5410 (
            .O(N__26141),
            .I(N__26106));
    Span12Mux_h I__5409 (
            .O(N__26138),
            .I(N__26101));
    Span12Mux_h I__5408 (
            .O(N__26133),
            .I(N__26101));
    LocalMux I__5407 (
            .O(N__26130),
            .I(N__26098));
    LocalMux I__5406 (
            .O(N__26127),
            .I(N__26095));
    Span4Mux_h I__5405 (
            .O(N__26124),
            .I(N__26090));
    Span4Mux_h I__5404 (
            .O(N__26121),
            .I(N__26090));
    Sp12to4 I__5403 (
            .O(N__26118),
            .I(N__26085));
    Sp12to4 I__5402 (
            .O(N__26113),
            .I(N__26085));
    Sp12to4 I__5401 (
            .O(N__26106),
            .I(N__26080));
    Span12Mux_v I__5400 (
            .O(N__26101),
            .I(N__26080));
    Span12Mux_h I__5399 (
            .O(N__26098),
            .I(N__26071));
    Span12Mux_h I__5398 (
            .O(N__26095),
            .I(N__26071));
    Sp12to4 I__5397 (
            .O(N__26090),
            .I(N__26071));
    Span12Mux_v I__5396 (
            .O(N__26085),
            .I(N__26071));
    Odrv12 I__5395 (
            .O(N__26080),
            .I(M_this_ppu_spr_addr_6));
    Odrv12 I__5394 (
            .O(N__26071),
            .I(M_this_ppu_spr_addr_6));
    InMux I__5393 (
            .O(N__26066),
            .I(N__26063));
    LocalMux I__5392 (
            .O(N__26063),
            .I(N__26060));
    Sp12to4 I__5391 (
            .O(N__26060),
            .I(N__26057));
    Span12Mux_v I__5390 (
            .O(N__26057),
            .I(N__26054));
    Odrv12 I__5389 (
            .O(N__26054),
            .I(\this_ppu.oam_cache.mem_0 ));
    InMux I__5388 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__5387 (
            .O(N__26048),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ));
    InMux I__5386 (
            .O(N__26045),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_0 ));
    InMux I__5385 (
            .O(N__26042),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_1 ));
    InMux I__5384 (
            .O(N__26039),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_2 ));
    InMux I__5383 (
            .O(N__26036),
            .I(\this_vga_signals.un1_M_vcounter_q_cry_3 ));
    InMux I__5382 (
            .O(N__26033),
            .I(N__26030));
    LocalMux I__5381 (
            .O(N__26030),
            .I(N__26027));
    Span4Mux_h I__5380 (
            .O(N__26027),
            .I(N__26024));
    Odrv4 I__5379 (
            .O(N__26024),
            .I(M_this_data_count_q_cry_3_THRU_CO));
    CascadeMux I__5378 (
            .O(N__26021),
            .I(N__26018));
    InMux I__5377 (
            .O(N__26018),
            .I(N__26015));
    LocalMux I__5376 (
            .O(N__26015),
            .I(N__26010));
    InMux I__5375 (
            .O(N__26014),
            .I(N__26005));
    InMux I__5374 (
            .O(N__26013),
            .I(N__26005));
    Odrv4 I__5373 (
            .O(N__26010),
            .I(M_this_data_count_qZ0Z_4));
    LocalMux I__5372 (
            .O(N__26005),
            .I(M_this_data_count_qZ0Z_4));
    CascadeMux I__5371 (
            .O(N__26000),
            .I(N__25997));
    InMux I__5370 (
            .O(N__25997),
            .I(N__25994));
    LocalMux I__5369 (
            .O(N__25994),
            .I(N__25991));
    Odrv12 I__5368 (
            .O(N__25991),
            .I(M_this_data_count_q_cry_4_THRU_CO));
    InMux I__5367 (
            .O(N__25988),
            .I(N__25985));
    LocalMux I__5366 (
            .O(N__25985),
            .I(N__25980));
    InMux I__5365 (
            .O(N__25984),
            .I(N__25975));
    InMux I__5364 (
            .O(N__25983),
            .I(N__25975));
    Odrv4 I__5363 (
            .O(N__25980),
            .I(M_this_data_count_qZ0Z_5));
    LocalMux I__5362 (
            .O(N__25975),
            .I(M_this_data_count_qZ0Z_5));
    InMux I__5361 (
            .O(N__25970),
            .I(N__25967));
    LocalMux I__5360 (
            .O(N__25967),
            .I(M_this_data_count_q_cry_8_THRU_CO));
    CascadeMux I__5359 (
            .O(N__25964),
            .I(N__25960));
    CascadeMux I__5358 (
            .O(N__25963),
            .I(N__25956));
    InMux I__5357 (
            .O(N__25960),
            .I(N__25953));
    InMux I__5356 (
            .O(N__25959),
            .I(N__25948));
    InMux I__5355 (
            .O(N__25956),
            .I(N__25948));
    LocalMux I__5354 (
            .O(N__25953),
            .I(M_this_data_count_qZ0Z_9));
    LocalMux I__5353 (
            .O(N__25948),
            .I(M_this_data_count_qZ0Z_9));
    InMux I__5352 (
            .O(N__25943),
            .I(N__25938));
    InMux I__5351 (
            .O(N__25942),
            .I(N__25933));
    InMux I__5350 (
            .O(N__25941),
            .I(N__25930));
    LocalMux I__5349 (
            .O(N__25938),
            .I(N__25927));
    InMux I__5348 (
            .O(N__25937),
            .I(N__25924));
    InMux I__5347 (
            .O(N__25936),
            .I(N__25921));
    LocalMux I__5346 (
            .O(N__25933),
            .I(\this_start_data_delay.M_last_qZ0 ));
    LocalMux I__5345 (
            .O(N__25930),
            .I(\this_start_data_delay.M_last_qZ0 ));
    Odrv4 I__5344 (
            .O(N__25927),
            .I(\this_start_data_delay.M_last_qZ0 ));
    LocalMux I__5343 (
            .O(N__25924),
            .I(\this_start_data_delay.M_last_qZ0 ));
    LocalMux I__5342 (
            .O(N__25921),
            .I(\this_start_data_delay.M_last_qZ0 ));
    CascadeMux I__5341 (
            .O(N__25910),
            .I(N_685_i_cascade_));
    CascadeMux I__5340 (
            .O(N__25907),
            .I(N__25904));
    InMux I__5339 (
            .O(N__25904),
            .I(N__25900));
    InMux I__5338 (
            .O(N__25903),
            .I(N__25896));
    LocalMux I__5337 (
            .O(N__25900),
            .I(N__25893));
    InMux I__5336 (
            .O(N__25899),
            .I(N__25890));
    LocalMux I__5335 (
            .O(N__25896),
            .I(M_this_data_count_qZ0Z_2));
    Odrv4 I__5334 (
            .O(N__25893),
            .I(M_this_data_count_qZ0Z_2));
    LocalMux I__5333 (
            .O(N__25890),
            .I(M_this_data_count_qZ0Z_2));
    InMux I__5332 (
            .O(N__25883),
            .I(N__25879));
    InMux I__5331 (
            .O(N__25882),
            .I(N__25875));
    LocalMux I__5330 (
            .O(N__25879),
            .I(N__25872));
    InMux I__5329 (
            .O(N__25878),
            .I(N__25869));
    LocalMux I__5328 (
            .O(N__25875),
            .I(M_this_data_count_qZ0Z_1));
    Odrv4 I__5327 (
            .O(N__25872),
            .I(M_this_data_count_qZ0Z_1));
    LocalMux I__5326 (
            .O(N__25869),
            .I(M_this_data_count_qZ0Z_1));
    InMux I__5325 (
            .O(N__25862),
            .I(N__25857));
    CascadeMux I__5324 (
            .O(N__25861),
            .I(N__25854));
    InMux I__5323 (
            .O(N__25860),
            .I(N__25851));
    LocalMux I__5322 (
            .O(N__25857),
            .I(N__25848));
    InMux I__5321 (
            .O(N__25854),
            .I(N__25845));
    LocalMux I__5320 (
            .O(N__25851),
            .I(M_this_data_count_qZ0Z_3));
    Odrv4 I__5319 (
            .O(N__25848),
            .I(M_this_data_count_qZ0Z_3));
    LocalMux I__5318 (
            .O(N__25845),
            .I(M_this_data_count_qZ0Z_3));
    InMux I__5317 (
            .O(N__25838),
            .I(N__25835));
    LocalMux I__5316 (
            .O(N__25835),
            .I(N__25830));
    InMux I__5315 (
            .O(N__25834),
            .I(N__25825));
    InMux I__5314 (
            .O(N__25833),
            .I(N__25825));
    Odrv4 I__5313 (
            .O(N__25830),
            .I(M_this_data_count_qZ0Z_0));
    LocalMux I__5312 (
            .O(N__25825),
            .I(M_this_data_count_qZ0Z_0));
    InMux I__5311 (
            .O(N__25820),
            .I(N__25817));
    LocalMux I__5310 (
            .O(N__25817),
            .I(\this_reset_cond.M_stage_qZ0Z_1 ));
    InMux I__5309 (
            .O(N__25814),
            .I(M_this_data_count_q_cry_8));
    InMux I__5308 (
            .O(N__25811),
            .I(M_this_data_count_q_cry_9));
    InMux I__5307 (
            .O(N__25808),
            .I(M_this_data_count_q_cry_10));
    IoInMux I__5306 (
            .O(N__25805),
            .I(N__25802));
    LocalMux I__5305 (
            .O(N__25802),
            .I(N__25792));
    SRMux I__5304 (
            .O(N__25801),
            .I(N__25789));
    SRMux I__5303 (
            .O(N__25800),
            .I(N__25784));
    SRMux I__5302 (
            .O(N__25799),
            .I(N__25781));
    SRMux I__5301 (
            .O(N__25798),
            .I(N__25778));
    SRMux I__5300 (
            .O(N__25797),
            .I(N__25773));
    SRMux I__5299 (
            .O(N__25796),
            .I(N__25770));
    SRMux I__5298 (
            .O(N__25795),
            .I(N__25767));
    IoSpan4Mux I__5297 (
            .O(N__25792),
            .I(N__25761));
    LocalMux I__5296 (
            .O(N__25789),
            .I(N__25758));
    SRMux I__5295 (
            .O(N__25788),
            .I(N__25755));
    SRMux I__5294 (
            .O(N__25787),
            .I(N__25752));
    LocalMux I__5293 (
            .O(N__25784),
            .I(N__25749));
    LocalMux I__5292 (
            .O(N__25781),
            .I(N__25744));
    LocalMux I__5291 (
            .O(N__25778),
            .I(N__25744));
    SRMux I__5290 (
            .O(N__25777),
            .I(N__25741));
    SRMux I__5289 (
            .O(N__25776),
            .I(N__25738));
    LocalMux I__5288 (
            .O(N__25773),
            .I(N__25733));
    LocalMux I__5287 (
            .O(N__25770),
            .I(N__25728));
    LocalMux I__5286 (
            .O(N__25767),
            .I(N__25728));
    SRMux I__5285 (
            .O(N__25766),
            .I(N__25725));
    SRMux I__5284 (
            .O(N__25765),
            .I(N__25714));
    SRMux I__5283 (
            .O(N__25764),
            .I(N__25711));
    Span4Mux_s3_h I__5282 (
            .O(N__25761),
            .I(N__25708));
    Span4Mux_s3_v I__5281 (
            .O(N__25758),
            .I(N__25701));
    LocalMux I__5280 (
            .O(N__25755),
            .I(N__25701));
    LocalMux I__5279 (
            .O(N__25752),
            .I(N__25701));
    Span4Mux_s3_v I__5278 (
            .O(N__25749),
            .I(N__25692));
    Span4Mux_s3_v I__5277 (
            .O(N__25744),
            .I(N__25692));
    LocalMux I__5276 (
            .O(N__25741),
            .I(N__25692));
    LocalMux I__5275 (
            .O(N__25738),
            .I(N__25692));
    SRMux I__5274 (
            .O(N__25737),
            .I(N__25689));
    SRMux I__5273 (
            .O(N__25736),
            .I(N__25686));
    Span4Mux_s3_v I__5272 (
            .O(N__25733),
            .I(N__25671));
    Span4Mux_s3_v I__5271 (
            .O(N__25728),
            .I(N__25671));
    LocalMux I__5270 (
            .O(N__25725),
            .I(N__25671));
    SRMux I__5269 (
            .O(N__25724),
            .I(N__25668));
    SRMux I__5268 (
            .O(N__25723),
            .I(N__25665));
    SRMux I__5267 (
            .O(N__25722),
            .I(N__25662));
    SRMux I__5266 (
            .O(N__25721),
            .I(N__25657));
    SRMux I__5265 (
            .O(N__25720),
            .I(N__25654));
    SRMux I__5264 (
            .O(N__25719),
            .I(N__25651));
    SRMux I__5263 (
            .O(N__25718),
            .I(N__25648));
    SRMux I__5262 (
            .O(N__25717),
            .I(N__25645));
    LocalMux I__5261 (
            .O(N__25714),
            .I(N__25640));
    LocalMux I__5260 (
            .O(N__25711),
            .I(N__25640));
    Span4Mux_h I__5259 (
            .O(N__25708),
            .I(N__25629));
    Span4Mux_v I__5258 (
            .O(N__25701),
            .I(N__25629));
    Span4Mux_v I__5257 (
            .O(N__25692),
            .I(N__25629));
    LocalMux I__5256 (
            .O(N__25689),
            .I(N__25629));
    LocalMux I__5255 (
            .O(N__25686),
            .I(N__25629));
    SRMux I__5254 (
            .O(N__25685),
            .I(N__25626));
    SRMux I__5253 (
            .O(N__25684),
            .I(N__25622));
    SRMux I__5252 (
            .O(N__25683),
            .I(N__25619));
    IoInMux I__5251 (
            .O(N__25682),
            .I(N__25615));
    SRMux I__5250 (
            .O(N__25681),
            .I(N__25612));
    SRMux I__5249 (
            .O(N__25680),
            .I(N__25609));
    SRMux I__5248 (
            .O(N__25679),
            .I(N__25606));
    SRMux I__5247 (
            .O(N__25678),
            .I(N__25603));
    Span4Mux_v I__5246 (
            .O(N__25671),
            .I(N__25594));
    LocalMux I__5245 (
            .O(N__25668),
            .I(N__25594));
    LocalMux I__5244 (
            .O(N__25665),
            .I(N__25589));
    LocalMux I__5243 (
            .O(N__25662),
            .I(N__25589));
    SRMux I__5242 (
            .O(N__25661),
            .I(N__25586));
    SRMux I__5241 (
            .O(N__25660),
            .I(N__25583));
    LocalMux I__5240 (
            .O(N__25657),
            .I(N__25575));
    LocalMux I__5239 (
            .O(N__25654),
            .I(N__25575));
    LocalMux I__5238 (
            .O(N__25651),
            .I(N__25570));
    LocalMux I__5237 (
            .O(N__25648),
            .I(N__25570));
    LocalMux I__5236 (
            .O(N__25645),
            .I(N__25567));
    Span4Mux_v I__5235 (
            .O(N__25640),
            .I(N__25560));
    Span4Mux_v I__5234 (
            .O(N__25629),
            .I(N__25560));
    LocalMux I__5233 (
            .O(N__25626),
            .I(N__25560));
    SRMux I__5232 (
            .O(N__25625),
            .I(N__25557));
    LocalMux I__5231 (
            .O(N__25622),
            .I(N__25554));
    LocalMux I__5230 (
            .O(N__25619),
            .I(N__25551));
    SRMux I__5229 (
            .O(N__25618),
            .I(N__25548));
    LocalMux I__5228 (
            .O(N__25615),
            .I(N__25545));
    LocalMux I__5227 (
            .O(N__25612),
            .I(N__25538));
    LocalMux I__5226 (
            .O(N__25609),
            .I(N__25538));
    LocalMux I__5225 (
            .O(N__25606),
            .I(N__25533));
    LocalMux I__5224 (
            .O(N__25603),
            .I(N__25533));
    SRMux I__5223 (
            .O(N__25602),
            .I(N__25530));
    SRMux I__5222 (
            .O(N__25601),
            .I(N__25527));
    SRMux I__5221 (
            .O(N__25600),
            .I(N__25524));
    SRMux I__5220 (
            .O(N__25599),
            .I(N__25521));
    Span4Mux_h I__5219 (
            .O(N__25594),
            .I(N__25516));
    Span4Mux_v I__5218 (
            .O(N__25589),
            .I(N__25516));
    LocalMux I__5217 (
            .O(N__25586),
            .I(N__25510));
    LocalMux I__5216 (
            .O(N__25583),
            .I(N__25510));
    SRMux I__5215 (
            .O(N__25582),
            .I(N__25507));
    SRMux I__5214 (
            .O(N__25581),
            .I(N__25504));
    SRMux I__5213 (
            .O(N__25580),
            .I(N__25500));
    Span4Mux_v I__5212 (
            .O(N__25575),
            .I(N__25497));
    Span4Mux_v I__5211 (
            .O(N__25570),
            .I(N__25494));
    Span4Mux_h I__5210 (
            .O(N__25567),
            .I(N__25487));
    Span4Mux_v I__5209 (
            .O(N__25560),
            .I(N__25487));
    LocalMux I__5208 (
            .O(N__25557),
            .I(N__25487));
    Span4Mux_v I__5207 (
            .O(N__25554),
            .I(N__25480));
    Span4Mux_v I__5206 (
            .O(N__25551),
            .I(N__25480));
    LocalMux I__5205 (
            .O(N__25548),
            .I(N__25480));
    IoSpan4Mux I__5204 (
            .O(N__25545),
            .I(N__25477));
    SRMux I__5203 (
            .O(N__25544),
            .I(N__25474));
    SRMux I__5202 (
            .O(N__25543),
            .I(N__25471));
    Span4Mux_v I__5201 (
            .O(N__25538),
            .I(N__25462));
    Span4Mux_v I__5200 (
            .O(N__25533),
            .I(N__25462));
    LocalMux I__5199 (
            .O(N__25530),
            .I(N__25462));
    LocalMux I__5198 (
            .O(N__25527),
            .I(N__25462));
    LocalMux I__5197 (
            .O(N__25524),
            .I(N__25457));
    LocalMux I__5196 (
            .O(N__25521),
            .I(N__25457));
    Span4Mux_v I__5195 (
            .O(N__25516),
            .I(N__25454));
    SRMux I__5194 (
            .O(N__25515),
            .I(N__25451));
    Span4Mux_v I__5193 (
            .O(N__25510),
            .I(N__25444));
    LocalMux I__5192 (
            .O(N__25507),
            .I(N__25444));
    LocalMux I__5191 (
            .O(N__25504),
            .I(N__25444));
    SRMux I__5190 (
            .O(N__25503),
            .I(N__25441));
    LocalMux I__5189 (
            .O(N__25500),
            .I(N__25438));
    Span4Mux_v I__5188 (
            .O(N__25497),
            .I(N__25431));
    Span4Mux_v I__5187 (
            .O(N__25494),
            .I(N__25431));
    Span4Mux_v I__5186 (
            .O(N__25487),
            .I(N__25431));
    Span4Mux_v I__5185 (
            .O(N__25480),
            .I(N__25428));
    Span4Mux_s3_h I__5184 (
            .O(N__25477),
            .I(N__25425));
    LocalMux I__5183 (
            .O(N__25474),
            .I(N__25420));
    LocalMux I__5182 (
            .O(N__25471),
            .I(N__25420));
    Span4Mux_v I__5181 (
            .O(N__25462),
            .I(N__25415));
    Span4Mux_v I__5180 (
            .O(N__25457),
            .I(N__25415));
    Span4Mux_v I__5179 (
            .O(N__25454),
            .I(N__25406));
    LocalMux I__5178 (
            .O(N__25451),
            .I(N__25406));
    Span4Mux_v I__5177 (
            .O(N__25444),
            .I(N__25406));
    LocalMux I__5176 (
            .O(N__25441),
            .I(N__25406));
    Span12Mux_h I__5175 (
            .O(N__25438),
            .I(N__25396));
    Span4Mux_h I__5174 (
            .O(N__25431),
            .I(N__25391));
    Span4Mux_h I__5173 (
            .O(N__25428),
            .I(N__25391));
    Span4Mux_h I__5172 (
            .O(N__25425),
            .I(N__25382));
    Span4Mux_v I__5171 (
            .O(N__25420),
            .I(N__25382));
    Span4Mux_v I__5170 (
            .O(N__25415),
            .I(N__25382));
    Span4Mux_v I__5169 (
            .O(N__25406),
            .I(N__25382));
    CascadeMux I__5168 (
            .O(N__25405),
            .I(N__25379));
    CascadeMux I__5167 (
            .O(N__25404),
            .I(N__25375));
    CascadeMux I__5166 (
            .O(N__25403),
            .I(N__25371));
    CascadeMux I__5165 (
            .O(N__25402),
            .I(N__25367));
    CascadeMux I__5164 (
            .O(N__25401),
            .I(N__25363));
    CascadeMux I__5163 (
            .O(N__25400),
            .I(N__25359));
    CascadeMux I__5162 (
            .O(N__25399),
            .I(N__25356));
    Span12Mux_v I__5161 (
            .O(N__25396),
            .I(N__25353));
    Span4Mux_h I__5160 (
            .O(N__25391),
            .I(N__25350));
    Span4Mux_h I__5159 (
            .O(N__25382),
            .I(N__25347));
    InMux I__5158 (
            .O(N__25379),
            .I(N__25332));
    InMux I__5157 (
            .O(N__25378),
            .I(N__25332));
    InMux I__5156 (
            .O(N__25375),
            .I(N__25332));
    InMux I__5155 (
            .O(N__25374),
            .I(N__25332));
    InMux I__5154 (
            .O(N__25371),
            .I(N__25332));
    InMux I__5153 (
            .O(N__25370),
            .I(N__25332));
    InMux I__5152 (
            .O(N__25367),
            .I(N__25332));
    InMux I__5151 (
            .O(N__25366),
            .I(N__25321));
    InMux I__5150 (
            .O(N__25363),
            .I(N__25321));
    InMux I__5149 (
            .O(N__25362),
            .I(N__25321));
    InMux I__5148 (
            .O(N__25359),
            .I(N__25321));
    InMux I__5147 (
            .O(N__25356),
            .I(N__25321));
    Odrv12 I__5146 (
            .O(N__25353),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5145 (
            .O(N__25350),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5144 (
            .O(N__25347),
            .I(CONSTANT_ONE_NET));
    LocalMux I__5143 (
            .O(N__25332),
            .I(CONSTANT_ONE_NET));
    LocalMux I__5142 (
            .O(N__25321),
            .I(CONSTANT_ONE_NET));
    InMux I__5141 (
            .O(N__25310),
            .I(M_this_data_count_q_cry_11));
    InMux I__5140 (
            .O(N__25307),
            .I(M_this_data_count_q_cry_12));
    CascadeMux I__5139 (
            .O(N__25304),
            .I(N__25301));
    InMux I__5138 (
            .O(N__25301),
            .I(N__25297));
    CascadeMux I__5137 (
            .O(N__25300),
            .I(N__25293));
    LocalMux I__5136 (
            .O(N__25297),
            .I(N__25288));
    InMux I__5135 (
            .O(N__25296),
            .I(N__25285));
    InMux I__5134 (
            .O(N__25293),
            .I(N__25278));
    InMux I__5133 (
            .O(N__25292),
            .I(N__25278));
    InMux I__5132 (
            .O(N__25291),
            .I(N__25278));
    Span4Mux_v I__5131 (
            .O(N__25288),
            .I(N__25275));
    LocalMux I__5130 (
            .O(N__25285),
            .I(N__25270));
    LocalMux I__5129 (
            .O(N__25278),
            .I(N__25270));
    Span4Mux_v I__5128 (
            .O(N__25275),
            .I(N__25267));
    Span4Mux_v I__5127 (
            .O(N__25270),
            .I(N__25264));
    Sp12to4 I__5126 (
            .O(N__25267),
            .I(N__25259));
    Sp12to4 I__5125 (
            .O(N__25264),
            .I(N__25259));
    Span12Mux_h I__5124 (
            .O(N__25259),
            .I(N__25256));
    Odrv12 I__5123 (
            .O(N__25256),
            .I(port_enb_c));
    InMux I__5122 (
            .O(N__25253),
            .I(N__25250));
    LocalMux I__5121 (
            .O(N__25250),
            .I(N__25243));
    InMux I__5120 (
            .O(N__25249),
            .I(N__25236));
    InMux I__5119 (
            .O(N__25248),
            .I(N__25236));
    InMux I__5118 (
            .O(N__25247),
            .I(N__25236));
    InMux I__5117 (
            .O(N__25246),
            .I(N__25233));
    Odrv4 I__5116 (
            .O(N__25243),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5115 (
            .O(N__25236),
            .I(M_this_delay_clk_out_0));
    LocalMux I__5114 (
            .O(N__25233),
            .I(M_this_delay_clk_out_0));
    InMux I__5113 (
            .O(N__25226),
            .I(N__25223));
    LocalMux I__5112 (
            .O(N__25223),
            .I(N__25220));
    Odrv4 I__5111 (
            .O(N__25220),
            .I(M_this_data_count_q_s_8));
    CascadeMux I__5110 (
            .O(N__25217),
            .I(N__25213));
    CascadeMux I__5109 (
            .O(N__25216),
            .I(N__25206));
    InMux I__5108 (
            .O(N__25213),
            .I(N__25201));
    InMux I__5107 (
            .O(N__25212),
            .I(N__25201));
    CascadeMux I__5106 (
            .O(N__25211),
            .I(N__25195));
    InMux I__5105 (
            .O(N__25210),
            .I(N__25190));
    InMux I__5104 (
            .O(N__25209),
            .I(N__25190));
    InMux I__5103 (
            .O(N__25206),
            .I(N__25187));
    LocalMux I__5102 (
            .O(N__25201),
            .I(N__25184));
    InMux I__5101 (
            .O(N__25200),
            .I(N__25179));
    InMux I__5100 (
            .O(N__25199),
            .I(N__25179));
    CascadeMux I__5099 (
            .O(N__25198),
            .I(N__25176));
    InMux I__5098 (
            .O(N__25195),
            .I(N__25173));
    LocalMux I__5097 (
            .O(N__25190),
            .I(N__25166));
    LocalMux I__5096 (
            .O(N__25187),
            .I(N__25166));
    Span4Mux_h I__5095 (
            .O(N__25184),
            .I(N__25166));
    LocalMux I__5094 (
            .O(N__25179),
            .I(N__25163));
    InMux I__5093 (
            .O(N__25176),
            .I(N__25160));
    LocalMux I__5092 (
            .O(N__25173),
            .I(N__25157));
    Span4Mux_v I__5091 (
            .O(N__25166),
            .I(N__25154));
    Span4Mux_v I__5090 (
            .O(N__25163),
            .I(N__25149));
    LocalMux I__5089 (
            .O(N__25160),
            .I(N__25149));
    Odrv4 I__5088 (
            .O(N__25157),
            .I(N_92));
    Odrv4 I__5087 (
            .O(N__25154),
            .I(N_92));
    Odrv4 I__5086 (
            .O(N__25149),
            .I(N_92));
    InMux I__5085 (
            .O(N__25142),
            .I(N__25138));
    InMux I__5084 (
            .O(N__25141),
            .I(N__25135));
    LocalMux I__5083 (
            .O(N__25138),
            .I(M_this_data_count_qZ0Z_8));
    LocalMux I__5082 (
            .O(N__25135),
            .I(M_this_data_count_qZ0Z_8));
    InMux I__5081 (
            .O(N__25130),
            .I(N__25127));
    LocalMux I__5080 (
            .O(N__25127),
            .I(N__25124));
    Span4Mux_h I__5079 (
            .O(N__25124),
            .I(N__25121));
    Odrv4 I__5078 (
            .O(N__25121),
            .I(M_this_data_count_q_cry_0_THRU_CO));
    InMux I__5077 (
            .O(N__25118),
            .I(M_this_data_count_q_cry_0));
    InMux I__5076 (
            .O(N__25115),
            .I(N__25112));
    LocalMux I__5075 (
            .O(N__25112),
            .I(N__25109));
    Odrv4 I__5074 (
            .O(N__25109),
            .I(M_this_data_count_q_cry_1_THRU_CO));
    InMux I__5073 (
            .O(N__25106),
            .I(M_this_data_count_q_cry_1));
    InMux I__5072 (
            .O(N__25103),
            .I(N__25100));
    LocalMux I__5071 (
            .O(N__25100),
            .I(N__25097));
    Odrv4 I__5070 (
            .O(N__25097),
            .I(M_this_data_count_q_cry_2_THRU_CO));
    InMux I__5069 (
            .O(N__25094),
            .I(M_this_data_count_q_cry_2));
    InMux I__5068 (
            .O(N__25091),
            .I(M_this_data_count_q_cry_3));
    InMux I__5067 (
            .O(N__25088),
            .I(M_this_data_count_q_cry_4));
    InMux I__5066 (
            .O(N__25085),
            .I(M_this_data_count_q_cry_5));
    CascadeMux I__5065 (
            .O(N__25082),
            .I(N__25079));
    InMux I__5064 (
            .O(N__25079),
            .I(N__25076));
    LocalMux I__5063 (
            .O(N__25076),
            .I(N__25073));
    Odrv4 I__5062 (
            .O(N__25073),
            .I(M_this_data_count_q_cry_6_THRU_CO));
    InMux I__5061 (
            .O(N__25070),
            .I(M_this_data_count_q_cry_6));
    InMux I__5060 (
            .O(N__25067),
            .I(bfn_15_20_0_));
    CascadeMux I__5059 (
            .O(N__25064),
            .I(N__25061));
    CascadeBuf I__5058 (
            .O(N__25061),
            .I(N__25058));
    CascadeMux I__5057 (
            .O(N__25058),
            .I(N__25055));
    InMux I__5056 (
            .O(N__25055),
            .I(N__25052));
    LocalMux I__5055 (
            .O(N__25052),
            .I(N__25049));
    Span4Mux_v I__5054 (
            .O(N__25049),
            .I(N__25046));
    Sp12to4 I__5053 (
            .O(N__25046),
            .I(N__25041));
    InMux I__5052 (
            .O(N__25045),
            .I(N__25038));
    InMux I__5051 (
            .O(N__25044),
            .I(N__25035));
    Span12Mux_h I__5050 (
            .O(N__25041),
            .I(N__25032));
    LocalMux I__5049 (
            .O(N__25038),
            .I(M_this_ppu_map_addr_4));
    LocalMux I__5048 (
            .O(N__25035),
            .I(M_this_ppu_map_addr_4));
    Odrv12 I__5047 (
            .O(N__25032),
            .I(M_this_ppu_map_addr_4));
    CascadeMux I__5046 (
            .O(N__25025),
            .I(N__25022));
    InMux I__5045 (
            .O(N__25022),
            .I(N__25019));
    LocalMux I__5044 (
            .O(N__25019),
            .I(N__25016));
    Odrv4 I__5043 (
            .O(N__25016),
            .I(\this_ppu.M_oam_cache_read_data_15 ));
    InMux I__5042 (
            .O(N__25013),
            .I(\this_ppu.offset_x_cry_6 ));
    InMux I__5041 (
            .O(N__25010),
            .I(N__25007));
    LocalMux I__5040 (
            .O(N__25007),
            .I(\this_ppu.offset_x_7 ));
    CascadeMux I__5039 (
            .O(N__25004),
            .I(N__25001));
    InMux I__5038 (
            .O(N__25001),
            .I(N__24998));
    LocalMux I__5037 (
            .O(N__24998),
            .I(M_this_scroll_qZ0Z_0));
    CascadeMux I__5036 (
            .O(N__24995),
            .I(N__24992));
    InMux I__5035 (
            .O(N__24992),
            .I(N__24989));
    LocalMux I__5034 (
            .O(N__24989),
            .I(M_this_scroll_qZ0Z_1));
    CascadeMux I__5033 (
            .O(N__24986),
            .I(N__24983));
    InMux I__5032 (
            .O(N__24983),
            .I(N__24980));
    LocalMux I__5031 (
            .O(N__24980),
            .I(M_this_scroll_qZ0Z_2));
    CascadeMux I__5030 (
            .O(N__24977),
            .I(N__24974));
    InMux I__5029 (
            .O(N__24974),
            .I(N__24971));
    LocalMux I__5028 (
            .O(N__24971),
            .I(N__24968));
    Odrv12 I__5027 (
            .O(N__24968),
            .I(M_this_scroll_qZ0Z_3));
    CascadeMux I__5026 (
            .O(N__24965),
            .I(N__24962));
    InMux I__5025 (
            .O(N__24962),
            .I(N__24959));
    LocalMux I__5024 (
            .O(N__24959),
            .I(M_this_scroll_qZ0Z_4));
    CascadeMux I__5023 (
            .O(N__24956),
            .I(N__24953));
    InMux I__5022 (
            .O(N__24953),
            .I(N__24950));
    LocalMux I__5021 (
            .O(N__24950),
            .I(M_this_scroll_qZ0Z_5));
    CascadeMux I__5020 (
            .O(N__24947),
            .I(N__24944));
    InMux I__5019 (
            .O(N__24944),
            .I(N__24941));
    LocalMux I__5018 (
            .O(N__24941),
            .I(M_this_scroll_qZ0Z_6));
    InMux I__5017 (
            .O(N__24938),
            .I(N__24935));
    LocalMux I__5016 (
            .O(N__24935),
            .I(M_this_scroll_qZ0Z_7));
    CascadeMux I__5015 (
            .O(N__24932),
            .I(\this_vga_signals.M_vcounter_d7lt8_0_cascade_ ));
    CascadeMux I__5014 (
            .O(N__24929),
            .I(N__24924));
    InMux I__5013 (
            .O(N__24928),
            .I(N__24919));
    InMux I__5012 (
            .O(N__24927),
            .I(N__24919));
    InMux I__5011 (
            .O(N__24924),
            .I(N__24916));
    LocalMux I__5010 (
            .O(N__24919),
            .I(N__24909));
    LocalMux I__5009 (
            .O(N__24916),
            .I(N__24906));
    InMux I__5008 (
            .O(N__24915),
            .I(N__24901));
    InMux I__5007 (
            .O(N__24914),
            .I(N__24901));
    InMux I__5006 (
            .O(N__24913),
            .I(N__24896));
    InMux I__5005 (
            .O(N__24912),
            .I(N__24896));
    Span4Mux_v I__5004 (
            .O(N__24909),
            .I(N__24891));
    Span4Mux_h I__5003 (
            .O(N__24906),
            .I(N__24891));
    LocalMux I__5002 (
            .O(N__24901),
            .I(\this_ppu.offset_x ));
    LocalMux I__5001 (
            .O(N__24896),
            .I(\this_ppu.offset_x ));
    Odrv4 I__5000 (
            .O(N__24891),
            .I(\this_ppu.offset_x ));
    InMux I__4999 (
            .O(N__24884),
            .I(N__24881));
    LocalMux I__4998 (
            .O(N__24881),
            .I(\this_ppu.M_oam_cache_read_data_i_8 ));
    InMux I__4997 (
            .O(N__24878),
            .I(N__24875));
    LocalMux I__4996 (
            .O(N__24875),
            .I(N__24872));
    Span4Mux_h I__4995 (
            .O(N__24872),
            .I(N__24869));
    Odrv4 I__4994 (
            .O(N__24869),
            .I(\this_ppu.M_oam_cache_read_data_i_9 ));
    CascadeMux I__4993 (
            .O(N__24866),
            .I(N__24859));
    InMux I__4992 (
            .O(N__24865),
            .I(N__24856));
    InMux I__4991 (
            .O(N__24864),
            .I(N__24853));
    InMux I__4990 (
            .O(N__24863),
            .I(N__24848));
    InMux I__4989 (
            .O(N__24862),
            .I(N__24848));
    InMux I__4988 (
            .O(N__24859),
            .I(N__24845));
    LocalMux I__4987 (
            .O(N__24856),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    LocalMux I__4986 (
            .O(N__24853),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    LocalMux I__4985 (
            .O(N__24848),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    LocalMux I__4984 (
            .O(N__24845),
            .I(\this_ppu.M_surface_x_qZ0Z_1 ));
    CascadeMux I__4983 (
            .O(N__24836),
            .I(N__24833));
    InMux I__4982 (
            .O(N__24833),
            .I(N__24829));
    CascadeMux I__4981 (
            .O(N__24832),
            .I(N__24826));
    LocalMux I__4980 (
            .O(N__24829),
            .I(N__24822));
    InMux I__4979 (
            .O(N__24826),
            .I(N__24819));
    CascadeMux I__4978 (
            .O(N__24825),
            .I(N__24816));
    Span4Mux_h I__4977 (
            .O(N__24822),
            .I(N__24809));
    LocalMux I__4976 (
            .O(N__24819),
            .I(N__24809));
    InMux I__4975 (
            .O(N__24816),
            .I(N__24806));
    CascadeMux I__4974 (
            .O(N__24815),
            .I(N__24803));
    CascadeMux I__4973 (
            .O(N__24814),
            .I(N__24798));
    Span4Mux_v I__4972 (
            .O(N__24809),
            .I(N__24791));
    LocalMux I__4971 (
            .O(N__24806),
            .I(N__24791));
    InMux I__4970 (
            .O(N__24803),
            .I(N__24788));
    CascadeMux I__4969 (
            .O(N__24802),
            .I(N__24785));
    CascadeMux I__4968 (
            .O(N__24801),
            .I(N__24781));
    InMux I__4967 (
            .O(N__24798),
            .I(N__24777));
    CascadeMux I__4966 (
            .O(N__24797),
            .I(N__24774));
    CascadeMux I__4965 (
            .O(N__24796),
            .I(N__24771));
    Span4Mux_v I__4964 (
            .O(N__24791),
            .I(N__24765));
    LocalMux I__4963 (
            .O(N__24788),
            .I(N__24765));
    InMux I__4962 (
            .O(N__24785),
            .I(N__24762));
    CascadeMux I__4961 (
            .O(N__24784),
            .I(N__24759));
    InMux I__4960 (
            .O(N__24781),
            .I(N__24755));
    CascadeMux I__4959 (
            .O(N__24780),
            .I(N__24752));
    LocalMux I__4958 (
            .O(N__24777),
            .I(N__24749));
    InMux I__4957 (
            .O(N__24774),
            .I(N__24746));
    InMux I__4956 (
            .O(N__24771),
            .I(N__24743));
    CascadeMux I__4955 (
            .O(N__24770),
            .I(N__24740));
    Span4Mux_h I__4954 (
            .O(N__24765),
            .I(N__24733));
    LocalMux I__4953 (
            .O(N__24762),
            .I(N__24733));
    InMux I__4952 (
            .O(N__24759),
            .I(N__24730));
    CascadeMux I__4951 (
            .O(N__24758),
            .I(N__24727));
    LocalMux I__4950 (
            .O(N__24755),
            .I(N__24724));
    InMux I__4949 (
            .O(N__24752),
            .I(N__24721));
    Span4Mux_h I__4948 (
            .O(N__24749),
            .I(N__24718));
    LocalMux I__4947 (
            .O(N__24746),
            .I(N__24715));
    LocalMux I__4946 (
            .O(N__24743),
            .I(N__24712));
    InMux I__4945 (
            .O(N__24740),
            .I(N__24709));
    CascadeMux I__4944 (
            .O(N__24739),
            .I(N__24706));
    CascadeMux I__4943 (
            .O(N__24738),
            .I(N__24703));
    Span4Mux_v I__4942 (
            .O(N__24733),
            .I(N__24698));
    LocalMux I__4941 (
            .O(N__24730),
            .I(N__24698));
    InMux I__4940 (
            .O(N__24727),
            .I(N__24695));
    Span4Mux_h I__4939 (
            .O(N__24724),
            .I(N__24691));
    LocalMux I__4938 (
            .O(N__24721),
            .I(N__24688));
    Span4Mux_v I__4937 (
            .O(N__24718),
            .I(N__24683));
    Span4Mux_h I__4936 (
            .O(N__24715),
            .I(N__24683));
    Span4Mux_h I__4935 (
            .O(N__24712),
            .I(N__24680));
    LocalMux I__4934 (
            .O(N__24709),
            .I(N__24677));
    InMux I__4933 (
            .O(N__24706),
            .I(N__24674));
    InMux I__4932 (
            .O(N__24703),
            .I(N__24671));
    Span4Mux_h I__4931 (
            .O(N__24698),
            .I(N__24666));
    LocalMux I__4930 (
            .O(N__24695),
            .I(N__24666));
    CascadeMux I__4929 (
            .O(N__24694),
            .I(N__24663));
    Span4Mux_h I__4928 (
            .O(N__24691),
            .I(N__24660));
    Span4Mux_h I__4927 (
            .O(N__24688),
            .I(N__24657));
    Span4Mux_v I__4926 (
            .O(N__24683),
            .I(N__24654));
    Span4Mux_v I__4925 (
            .O(N__24680),
            .I(N__24649));
    Span4Mux_h I__4924 (
            .O(N__24677),
            .I(N__24649));
    LocalMux I__4923 (
            .O(N__24674),
            .I(N__24646));
    LocalMux I__4922 (
            .O(N__24671),
            .I(N__24643));
    Span4Mux_v I__4921 (
            .O(N__24666),
            .I(N__24640));
    InMux I__4920 (
            .O(N__24663),
            .I(N__24637));
    Sp12to4 I__4919 (
            .O(N__24660),
            .I(N__24634));
    Span4Mux_h I__4918 (
            .O(N__24657),
            .I(N__24631));
    Span4Mux_v I__4917 (
            .O(N__24654),
            .I(N__24628));
    Span4Mux_h I__4916 (
            .O(N__24649),
            .I(N__24625));
    Span12Mux_s10_h I__4915 (
            .O(N__24646),
            .I(N__24622));
    Span12Mux_s9_h I__4914 (
            .O(N__24643),
            .I(N__24619));
    Sp12to4 I__4913 (
            .O(N__24640),
            .I(N__24614));
    LocalMux I__4912 (
            .O(N__24637),
            .I(N__24614));
    Span12Mux_v I__4911 (
            .O(N__24634),
            .I(N__24609));
    Sp12to4 I__4910 (
            .O(N__24631),
            .I(N__24609));
    Span4Mux_h I__4909 (
            .O(N__24628),
            .I(N__24604));
    Span4Mux_v I__4908 (
            .O(N__24625),
            .I(N__24604));
    Span12Mux_v I__4907 (
            .O(N__24622),
            .I(N__24597));
    Span12Mux_v I__4906 (
            .O(N__24619),
            .I(N__24597));
    Span12Mux_s10_h I__4905 (
            .O(N__24614),
            .I(N__24597));
    Odrv12 I__4904 (
            .O(N__24609),
            .I(M_this_ppu_spr_addr_1));
    Odrv4 I__4903 (
            .O(N__24604),
            .I(M_this_ppu_spr_addr_1));
    Odrv12 I__4902 (
            .O(N__24597),
            .I(M_this_ppu_spr_addr_1));
    InMux I__4901 (
            .O(N__24590),
            .I(\this_ppu.offset_x_cry_0 ));
    InMux I__4900 (
            .O(N__24587),
            .I(N__24584));
    LocalMux I__4899 (
            .O(N__24584),
            .I(N__24581));
    Odrv12 I__4898 (
            .O(N__24581),
            .I(\this_ppu.M_oam_cache_read_data_i_10 ));
    CascadeMux I__4897 (
            .O(N__24578),
            .I(N__24575));
    InMux I__4896 (
            .O(N__24575),
            .I(N__24568));
    InMux I__4895 (
            .O(N__24574),
            .I(N__24565));
    InMux I__4894 (
            .O(N__24573),
            .I(N__24558));
    InMux I__4893 (
            .O(N__24572),
            .I(N__24558));
    InMux I__4892 (
            .O(N__24571),
            .I(N__24558));
    LocalMux I__4891 (
            .O(N__24568),
            .I(N__24555));
    LocalMux I__4890 (
            .O(N__24565),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    LocalMux I__4889 (
            .O(N__24558),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    Odrv4 I__4888 (
            .O(N__24555),
            .I(\this_ppu.M_surface_x_qZ0Z_2 ));
    CascadeMux I__4887 (
            .O(N__24548),
            .I(N__24545));
    InMux I__4886 (
            .O(N__24545),
            .I(N__24541));
    CascadeMux I__4885 (
            .O(N__24544),
            .I(N__24538));
    LocalMux I__4884 (
            .O(N__24541),
            .I(N__24533));
    InMux I__4883 (
            .O(N__24538),
            .I(N__24530));
    CascadeMux I__4882 (
            .O(N__24537),
            .I(N__24527));
    CascadeMux I__4881 (
            .O(N__24536),
            .I(N__24522));
    Span4Mux_v I__4880 (
            .O(N__24533),
            .I(N__24517));
    LocalMux I__4879 (
            .O(N__24530),
            .I(N__24517));
    InMux I__4878 (
            .O(N__24527),
            .I(N__24514));
    CascadeMux I__4877 (
            .O(N__24526),
            .I(N__24511));
    CascadeMux I__4876 (
            .O(N__24525),
            .I(N__24507));
    InMux I__4875 (
            .O(N__24522),
            .I(N__24503));
    Span4Mux_h I__4874 (
            .O(N__24517),
            .I(N__24496));
    LocalMux I__4873 (
            .O(N__24514),
            .I(N__24496));
    InMux I__4872 (
            .O(N__24511),
            .I(N__24493));
    CascadeMux I__4871 (
            .O(N__24510),
            .I(N__24490));
    InMux I__4870 (
            .O(N__24507),
            .I(N__24487));
    CascadeMux I__4869 (
            .O(N__24506),
            .I(N__24484));
    LocalMux I__4868 (
            .O(N__24503),
            .I(N__24477));
    CascadeMux I__4867 (
            .O(N__24502),
            .I(N__24474));
    CascadeMux I__4866 (
            .O(N__24501),
            .I(N__24471));
    Span4Mux_v I__4865 (
            .O(N__24496),
            .I(N__24466));
    LocalMux I__4864 (
            .O(N__24493),
            .I(N__24466));
    InMux I__4863 (
            .O(N__24490),
            .I(N__24463));
    LocalMux I__4862 (
            .O(N__24487),
            .I(N__24459));
    InMux I__4861 (
            .O(N__24484),
            .I(N__24456));
    CascadeMux I__4860 (
            .O(N__24483),
            .I(N__24453));
    CascadeMux I__4859 (
            .O(N__24482),
            .I(N__24450));
    CascadeMux I__4858 (
            .O(N__24481),
            .I(N__24447));
    CascadeMux I__4857 (
            .O(N__24480),
            .I(N__24444));
    Span4Mux_s2_v I__4856 (
            .O(N__24477),
            .I(N__24440));
    InMux I__4855 (
            .O(N__24474),
            .I(N__24437));
    InMux I__4854 (
            .O(N__24471),
            .I(N__24434));
    Span4Mux_h I__4853 (
            .O(N__24466),
            .I(N__24429));
    LocalMux I__4852 (
            .O(N__24463),
            .I(N__24429));
    CascadeMux I__4851 (
            .O(N__24462),
            .I(N__24426));
    Span4Mux_s0_v I__4850 (
            .O(N__24459),
            .I(N__24423));
    LocalMux I__4849 (
            .O(N__24456),
            .I(N__24420));
    InMux I__4848 (
            .O(N__24453),
            .I(N__24417));
    InMux I__4847 (
            .O(N__24450),
            .I(N__24414));
    InMux I__4846 (
            .O(N__24447),
            .I(N__24411));
    InMux I__4845 (
            .O(N__24444),
            .I(N__24408));
    CascadeMux I__4844 (
            .O(N__24443),
            .I(N__24405));
    Sp12to4 I__4843 (
            .O(N__24440),
            .I(N__24400));
    LocalMux I__4842 (
            .O(N__24437),
            .I(N__24400));
    LocalMux I__4841 (
            .O(N__24434),
            .I(N__24397));
    Span4Mux_v I__4840 (
            .O(N__24429),
            .I(N__24394));
    InMux I__4839 (
            .O(N__24426),
            .I(N__24391));
    Span4Mux_v I__4838 (
            .O(N__24423),
            .I(N__24384));
    Span4Mux_h I__4837 (
            .O(N__24420),
            .I(N__24384));
    LocalMux I__4836 (
            .O(N__24417),
            .I(N__24384));
    LocalMux I__4835 (
            .O(N__24414),
            .I(N__24381));
    LocalMux I__4834 (
            .O(N__24411),
            .I(N__24378));
    LocalMux I__4833 (
            .O(N__24408),
            .I(N__24375));
    InMux I__4832 (
            .O(N__24405),
            .I(N__24372));
    Span12Mux_h I__4831 (
            .O(N__24400),
            .I(N__24367));
    Span12Mux_h I__4830 (
            .O(N__24397),
            .I(N__24367));
    Sp12to4 I__4829 (
            .O(N__24394),
            .I(N__24362));
    LocalMux I__4828 (
            .O(N__24391),
            .I(N__24362));
    Sp12to4 I__4827 (
            .O(N__24384),
            .I(N__24359));
    Sp12to4 I__4826 (
            .O(N__24381),
            .I(N__24352));
    Sp12to4 I__4825 (
            .O(N__24378),
            .I(N__24352));
    Sp12to4 I__4824 (
            .O(N__24375),
            .I(N__24352));
    LocalMux I__4823 (
            .O(N__24372),
            .I(N__24349));
    Span12Mux_v I__4822 (
            .O(N__24367),
            .I(N__24344));
    Span12Mux_h I__4821 (
            .O(N__24362),
            .I(N__24344));
    Span12Mux_v I__4820 (
            .O(N__24359),
            .I(N__24337));
    Span12Mux_v I__4819 (
            .O(N__24352),
            .I(N__24337));
    Span12Mux_s11_h I__4818 (
            .O(N__24349),
            .I(N__24337));
    Odrv12 I__4817 (
            .O(N__24344),
            .I(M_this_ppu_spr_addr_2));
    Odrv12 I__4816 (
            .O(N__24337),
            .I(M_this_ppu_spr_addr_2));
    InMux I__4815 (
            .O(N__24332),
            .I(\this_ppu.offset_x_cry_1 ));
    CascadeMux I__4814 (
            .O(N__24329),
            .I(N__24325));
    CascadeMux I__4813 (
            .O(N__24328),
            .I(N__24322));
    CascadeBuf I__4812 (
            .O(N__24325),
            .I(N__24319));
    InMux I__4811 (
            .O(N__24322),
            .I(N__24316));
    CascadeMux I__4810 (
            .O(N__24319),
            .I(N__24313));
    LocalMux I__4809 (
            .O(N__24316),
            .I(N__24310));
    InMux I__4808 (
            .O(N__24313),
            .I(N__24307));
    Span4Mux_v I__4807 (
            .O(N__24310),
            .I(N__24300));
    LocalMux I__4806 (
            .O(N__24307),
            .I(N__24297));
    InMux I__4805 (
            .O(N__24306),
            .I(N__24292));
    InMux I__4804 (
            .O(N__24305),
            .I(N__24292));
    InMux I__4803 (
            .O(N__24304),
            .I(N__24287));
    InMux I__4802 (
            .O(N__24303),
            .I(N__24287));
    Sp12to4 I__4801 (
            .O(N__24300),
            .I(N__24282));
    Span12Mux_v I__4800 (
            .O(N__24297),
            .I(N__24282));
    LocalMux I__4799 (
            .O(N__24292),
            .I(M_this_ppu_map_addr_0));
    LocalMux I__4798 (
            .O(N__24287),
            .I(M_this_ppu_map_addr_0));
    Odrv12 I__4797 (
            .O(N__24282),
            .I(M_this_ppu_map_addr_0));
    InMux I__4796 (
            .O(N__24275),
            .I(N__24272));
    LocalMux I__4795 (
            .O(N__24272),
            .I(\this_ppu.offset_x_3 ));
    InMux I__4794 (
            .O(N__24269),
            .I(\this_ppu.offset_x_cry_2 ));
    CascadeMux I__4793 (
            .O(N__24266),
            .I(N__24263));
    CascadeBuf I__4792 (
            .O(N__24263),
            .I(N__24260));
    CascadeMux I__4791 (
            .O(N__24260),
            .I(N__24257));
    InMux I__4790 (
            .O(N__24257),
            .I(N__24254));
    LocalMux I__4789 (
            .O(N__24254),
            .I(N__24249));
    CascadeMux I__4788 (
            .O(N__24253),
            .I(N__24246));
    CascadeMux I__4787 (
            .O(N__24252),
            .I(N__24240));
    Sp12to4 I__4786 (
            .O(N__24249),
            .I(N__24237));
    InMux I__4785 (
            .O(N__24246),
            .I(N__24234));
    InMux I__4784 (
            .O(N__24245),
            .I(N__24231));
    InMux I__4783 (
            .O(N__24244),
            .I(N__24226));
    InMux I__4782 (
            .O(N__24243),
            .I(N__24226));
    InMux I__4781 (
            .O(N__24240),
            .I(N__24223));
    Span12Mux_v I__4780 (
            .O(N__24237),
            .I(N__24220));
    LocalMux I__4779 (
            .O(N__24234),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4778 (
            .O(N__24231),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4777 (
            .O(N__24226),
            .I(M_this_ppu_map_addr_1));
    LocalMux I__4776 (
            .O(N__24223),
            .I(M_this_ppu_map_addr_1));
    Odrv12 I__4775 (
            .O(N__24220),
            .I(M_this_ppu_map_addr_1));
    InMux I__4774 (
            .O(N__24209),
            .I(N__24206));
    LocalMux I__4773 (
            .O(N__24206),
            .I(\this_ppu.offset_x_4 ));
    InMux I__4772 (
            .O(N__24203),
            .I(\this_ppu.offset_x_cry_3 ));
    InMux I__4771 (
            .O(N__24200),
            .I(N__24197));
    LocalMux I__4770 (
            .O(N__24197),
            .I(N__24194));
    Span4Mux_h I__4769 (
            .O(N__24194),
            .I(N__24191));
    Odrv4 I__4768 (
            .O(N__24191),
            .I(\this_ppu.M_oam_cache_read_data_i_13 ));
    CascadeMux I__4767 (
            .O(N__24188),
            .I(N__24185));
    CascadeBuf I__4766 (
            .O(N__24185),
            .I(N__24182));
    CascadeMux I__4765 (
            .O(N__24182),
            .I(N__24178));
    CascadeMux I__4764 (
            .O(N__24181),
            .I(N__24175));
    InMux I__4763 (
            .O(N__24178),
            .I(N__24172));
    InMux I__4762 (
            .O(N__24175),
            .I(N__24169));
    LocalMux I__4761 (
            .O(N__24172),
            .I(N__24166));
    LocalMux I__4760 (
            .O(N__24169),
            .I(N__24160));
    Span12Mux_s7_h I__4759 (
            .O(N__24166),
            .I(N__24157));
    InMux I__4758 (
            .O(N__24165),
            .I(N__24154));
    InMux I__4757 (
            .O(N__24164),
            .I(N__24151));
    InMux I__4756 (
            .O(N__24163),
            .I(N__24148));
    Span4Mux_h I__4755 (
            .O(N__24160),
            .I(N__24145));
    Span12Mux_h I__4754 (
            .O(N__24157),
            .I(N__24142));
    LocalMux I__4753 (
            .O(N__24154),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__4752 (
            .O(N__24151),
            .I(M_this_ppu_map_addr_2));
    LocalMux I__4751 (
            .O(N__24148),
            .I(M_this_ppu_map_addr_2));
    Odrv4 I__4750 (
            .O(N__24145),
            .I(M_this_ppu_map_addr_2));
    Odrv12 I__4749 (
            .O(N__24142),
            .I(M_this_ppu_map_addr_2));
    InMux I__4748 (
            .O(N__24131),
            .I(N__24128));
    LocalMux I__4747 (
            .O(N__24128),
            .I(\this_ppu.offset_x_5 ));
    InMux I__4746 (
            .O(N__24125),
            .I(\this_ppu.offset_x_cry_4 ));
    InMux I__4745 (
            .O(N__24122),
            .I(N__24119));
    LocalMux I__4744 (
            .O(N__24119),
            .I(N__24116));
    Span4Mux_v I__4743 (
            .O(N__24116),
            .I(N__24113));
    Odrv4 I__4742 (
            .O(N__24113),
            .I(\this_ppu.M_oam_cache_read_data_i_14 ));
    CascadeMux I__4741 (
            .O(N__24110),
            .I(N__24107));
    CascadeBuf I__4740 (
            .O(N__24107),
            .I(N__24104));
    CascadeMux I__4739 (
            .O(N__24104),
            .I(N__24100));
    CascadeMux I__4738 (
            .O(N__24103),
            .I(N__24097));
    InMux I__4737 (
            .O(N__24100),
            .I(N__24094));
    InMux I__4736 (
            .O(N__24097),
            .I(N__24090));
    LocalMux I__4735 (
            .O(N__24094),
            .I(N__24087));
    CascadeMux I__4734 (
            .O(N__24093),
            .I(N__24083));
    LocalMux I__4733 (
            .O(N__24090),
            .I(N__24080));
    Span12Mux_s7_v I__4732 (
            .O(N__24087),
            .I(N__24077));
    InMux I__4731 (
            .O(N__24086),
            .I(N__24072));
    InMux I__4730 (
            .O(N__24083),
            .I(N__24072));
    Span4Mux_h I__4729 (
            .O(N__24080),
            .I(N__24069));
    Span12Mux_h I__4728 (
            .O(N__24077),
            .I(N__24066));
    LocalMux I__4727 (
            .O(N__24072),
            .I(M_this_ppu_map_addr_3));
    Odrv4 I__4726 (
            .O(N__24069),
            .I(M_this_ppu_map_addr_3));
    Odrv12 I__4725 (
            .O(N__24066),
            .I(M_this_ppu_map_addr_3));
    InMux I__4724 (
            .O(N__24059),
            .I(N__24056));
    LocalMux I__4723 (
            .O(N__24056),
            .I(\this_ppu.offset_x_6 ));
    InMux I__4722 (
            .O(N__24053),
            .I(\this_ppu.offset_x_cry_5 ));
    InMux I__4721 (
            .O(N__24050),
            .I(N__24046));
    CascadeMux I__4720 (
            .O(N__24049),
            .I(N__24043));
    LocalMux I__4719 (
            .O(N__24046),
            .I(N__24040));
    InMux I__4718 (
            .O(N__24043),
            .I(N__24037));
    Span4Mux_v I__4717 (
            .O(N__24040),
            .I(N__24033));
    LocalMux I__4716 (
            .O(N__24037),
            .I(N__24030));
    InMux I__4715 (
            .O(N__24036),
            .I(N__24027));
    Span4Mux_h I__4714 (
            .O(N__24033),
            .I(N__24022));
    Span4Mux_v I__4713 (
            .O(N__24030),
            .I(N__24022));
    LocalMux I__4712 (
            .O(N__24027),
            .I(M_this_ctrl_flags_qZ0Z_6));
    Odrv4 I__4711 (
            .O(N__24022),
            .I(M_this_ctrl_flags_qZ0Z_6));
    InMux I__4710 (
            .O(N__24017),
            .I(N__24014));
    LocalMux I__4709 (
            .O(N__24014),
            .I(N__24011));
    Span12Mux_v I__4708 (
            .O(N__24011),
            .I(N__24008));
    Odrv12 I__4707 (
            .O(N__24008),
            .I(M_this_oam_ram_read_data_13));
    CEMux I__4706 (
            .O(N__24005),
            .I(N__24002));
    LocalMux I__4705 (
            .O(N__24002),
            .I(N__23984));
    InMux I__4704 (
            .O(N__24001),
            .I(N__23968));
    InMux I__4703 (
            .O(N__24000),
            .I(N__23959));
    InMux I__4702 (
            .O(N__23999),
            .I(N__23959));
    InMux I__4701 (
            .O(N__23998),
            .I(N__23959));
    InMux I__4700 (
            .O(N__23997),
            .I(N__23959));
    InMux I__4699 (
            .O(N__23996),
            .I(N__23956));
    InMux I__4698 (
            .O(N__23995),
            .I(N__23952));
    InMux I__4697 (
            .O(N__23994),
            .I(N__23935));
    InMux I__4696 (
            .O(N__23993),
            .I(N__23935));
    InMux I__4695 (
            .O(N__23992),
            .I(N__23935));
    InMux I__4694 (
            .O(N__23991),
            .I(N__23935));
    InMux I__4693 (
            .O(N__23990),
            .I(N__23935));
    InMux I__4692 (
            .O(N__23989),
            .I(N__23935));
    InMux I__4691 (
            .O(N__23988),
            .I(N__23935));
    InMux I__4690 (
            .O(N__23987),
            .I(N__23932));
    Span4Mux_v I__4689 (
            .O(N__23984),
            .I(N__23929));
    InMux I__4688 (
            .O(N__23983),
            .I(N__23924));
    InMux I__4687 (
            .O(N__23982),
            .I(N__23924));
    InMux I__4686 (
            .O(N__23981),
            .I(N__23913));
    InMux I__4685 (
            .O(N__23980),
            .I(N__23913));
    InMux I__4684 (
            .O(N__23979),
            .I(N__23913));
    InMux I__4683 (
            .O(N__23978),
            .I(N__23913));
    InMux I__4682 (
            .O(N__23977),
            .I(N__23913));
    InMux I__4681 (
            .O(N__23976),
            .I(N__23904));
    InMux I__4680 (
            .O(N__23975),
            .I(N__23904));
    InMux I__4679 (
            .O(N__23974),
            .I(N__23904));
    InMux I__4678 (
            .O(N__23973),
            .I(N__23904));
    InMux I__4677 (
            .O(N__23972),
            .I(N__23899));
    InMux I__4676 (
            .O(N__23971),
            .I(N__23899));
    LocalMux I__4675 (
            .O(N__23968),
            .I(N__23894));
    LocalMux I__4674 (
            .O(N__23959),
            .I(N__23894));
    LocalMux I__4673 (
            .O(N__23956),
            .I(N__23891));
    InMux I__4672 (
            .O(N__23955),
            .I(N__23888));
    LocalMux I__4671 (
            .O(N__23952),
            .I(N__23879));
    InMux I__4670 (
            .O(N__23951),
            .I(N__23876));
    CEMux I__4669 (
            .O(N__23950),
            .I(N__23873));
    LocalMux I__4668 (
            .O(N__23935),
            .I(N__23870));
    LocalMux I__4667 (
            .O(N__23932),
            .I(N__23867));
    Span4Mux_v I__4666 (
            .O(N__23929),
            .I(N__23860));
    LocalMux I__4665 (
            .O(N__23924),
            .I(N__23860));
    LocalMux I__4664 (
            .O(N__23913),
            .I(N__23860));
    LocalMux I__4663 (
            .O(N__23904),
            .I(N__23855));
    LocalMux I__4662 (
            .O(N__23899),
            .I(N__23855));
    Span4Mux_v I__4661 (
            .O(N__23894),
            .I(N__23850));
    Span4Mux_v I__4660 (
            .O(N__23891),
            .I(N__23850));
    LocalMux I__4659 (
            .O(N__23888),
            .I(N__23846));
    InMux I__4658 (
            .O(N__23887),
            .I(N__23839));
    InMux I__4657 (
            .O(N__23886),
            .I(N__23839));
    InMux I__4656 (
            .O(N__23885),
            .I(N__23839));
    InMux I__4655 (
            .O(N__23884),
            .I(N__23832));
    InMux I__4654 (
            .O(N__23883),
            .I(N__23832));
    InMux I__4653 (
            .O(N__23882),
            .I(N__23832));
    Span4Mux_v I__4652 (
            .O(N__23879),
            .I(N__23827));
    LocalMux I__4651 (
            .O(N__23876),
            .I(N__23827));
    LocalMux I__4650 (
            .O(N__23873),
            .I(N__23824));
    Span4Mux_v I__4649 (
            .O(N__23870),
            .I(N__23817));
    Span4Mux_h I__4648 (
            .O(N__23867),
            .I(N__23817));
    Span4Mux_v I__4647 (
            .O(N__23860),
            .I(N__23817));
    Span12Mux_s6_v I__4646 (
            .O(N__23855),
            .I(N__23814));
    Span4Mux_h I__4645 (
            .O(N__23850),
            .I(N__23811));
    InMux I__4644 (
            .O(N__23849),
            .I(N__23808));
    Span4Mux_h I__4643 (
            .O(N__23846),
            .I(N__23805));
    LocalMux I__4642 (
            .O(N__23839),
            .I(N__23798));
    LocalMux I__4641 (
            .O(N__23832),
            .I(N__23798));
    Span4Mux_h I__4640 (
            .O(N__23827),
            .I(N__23798));
    Odrv12 I__4639 (
            .O(N__23824),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4638 (
            .O(N__23817),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv12 I__4637 (
            .O(N__23814),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4636 (
            .O(N__23811),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    LocalMux I__4635 (
            .O(N__23808),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4634 (
            .O(N__23805),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    Odrv4 I__4633 (
            .O(N__23798),
            .I(\this_ppu.M_state_qZ0Z_3 ));
    InMux I__4632 (
            .O(N__23783),
            .I(N__23780));
    LocalMux I__4631 (
            .O(N__23780),
            .I(N__23777));
    Span4Mux_v I__4630 (
            .O(N__23777),
            .I(N__23774));
    Span4Mux_v I__4629 (
            .O(N__23774),
            .I(N__23771));
    Span4Mux_h I__4628 (
            .O(N__23771),
            .I(N__23768));
    Odrv4 I__4627 (
            .O(N__23768),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_13 ));
    CascadeMux I__4626 (
            .O(N__23765),
            .I(N__23760));
    InMux I__4625 (
            .O(N__23764),
            .I(N__23752));
    InMux I__4624 (
            .O(N__23763),
            .I(N__23752));
    InMux I__4623 (
            .O(N__23760),
            .I(N__23749));
    InMux I__4622 (
            .O(N__23759),
            .I(N__23746));
    InMux I__4621 (
            .O(N__23758),
            .I(N__23743));
    InMux I__4620 (
            .O(N__23757),
            .I(N__23740));
    LocalMux I__4619 (
            .O(N__23752),
            .I(N__23737));
    LocalMux I__4618 (
            .O(N__23749),
            .I(N__23734));
    LocalMux I__4617 (
            .O(N__23746),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__4616 (
            .O(N__23743),
            .I(M_this_oam_address_qZ0Z_1));
    LocalMux I__4615 (
            .O(N__23740),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__4614 (
            .O(N__23737),
            .I(M_this_oam_address_qZ0Z_1));
    Odrv4 I__4613 (
            .O(N__23734),
            .I(M_this_oam_address_qZ0Z_1));
    InMux I__4612 (
            .O(N__23723),
            .I(N__23716));
    InMux I__4611 (
            .O(N__23722),
            .I(N__23713));
    InMux I__4610 (
            .O(N__23721),
            .I(N__23710));
    InMux I__4609 (
            .O(N__23720),
            .I(N__23705));
    InMux I__4608 (
            .O(N__23719),
            .I(N__23705));
    LocalMux I__4607 (
            .O(N__23716),
            .I(N__23699));
    LocalMux I__4606 (
            .O(N__23713),
            .I(N__23699));
    LocalMux I__4605 (
            .O(N__23710),
            .I(N__23694));
    LocalMux I__4604 (
            .O(N__23705),
            .I(N__23694));
    InMux I__4603 (
            .O(N__23704),
            .I(N__23690));
    Span4Mux_h I__4602 (
            .O(N__23699),
            .I(N__23687));
    Span4Mux_v I__4601 (
            .O(N__23694),
            .I(N__23684));
    InMux I__4600 (
            .O(N__23693),
            .I(N__23681));
    LocalMux I__4599 (
            .O(N__23690),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__4598 (
            .O(N__23687),
            .I(M_this_oam_address_qZ0Z_0));
    Odrv4 I__4597 (
            .O(N__23684),
            .I(M_this_oam_address_qZ0Z_0));
    LocalMux I__4596 (
            .O(N__23681),
            .I(M_this_oam_address_qZ0Z_0));
    CascadeMux I__4595 (
            .O(N__23672),
            .I(N__23668));
    CascadeMux I__4594 (
            .O(N__23671),
            .I(N__23664));
    InMux I__4593 (
            .O(N__23668),
            .I(N__23659));
    InMux I__4592 (
            .O(N__23667),
            .I(N__23655));
    InMux I__4591 (
            .O(N__23664),
            .I(N__23652));
    InMux I__4590 (
            .O(N__23663),
            .I(N__23647));
    InMux I__4589 (
            .O(N__23662),
            .I(N__23647));
    LocalMux I__4588 (
            .O(N__23659),
            .I(N__23644));
    InMux I__4587 (
            .O(N__23658),
            .I(N__23641));
    LocalMux I__4586 (
            .O(N__23655),
            .I(N__23634));
    LocalMux I__4585 (
            .O(N__23652),
            .I(N__23634));
    LocalMux I__4584 (
            .O(N__23647),
            .I(N__23634));
    Span4Mux_v I__4583 (
            .O(N__23644),
            .I(N__23631));
    LocalMux I__4582 (
            .O(N__23641),
            .I(N__23626));
    Span4Mux_v I__4581 (
            .O(N__23634),
            .I(N__23626));
    Odrv4 I__4580 (
            .O(N__23631),
            .I(N_222_0));
    Odrv4 I__4579 (
            .O(N__23626),
            .I(N_222_0));
    CEMux I__4578 (
            .O(N__23621),
            .I(N__23616));
    CEMux I__4577 (
            .O(N__23620),
            .I(N__23613));
    CEMux I__4576 (
            .O(N__23619),
            .I(N__23610));
    LocalMux I__4575 (
            .O(N__23616),
            .I(N__23607));
    LocalMux I__4574 (
            .O(N__23613),
            .I(N__23603));
    LocalMux I__4573 (
            .O(N__23610),
            .I(N__23600));
    Span4Mux_v I__4572 (
            .O(N__23607),
            .I(N__23597));
    CEMux I__4571 (
            .O(N__23606),
            .I(N__23594));
    Span4Mux_v I__4570 (
            .O(N__23603),
            .I(N__23589));
    Span4Mux_v I__4569 (
            .O(N__23600),
            .I(N__23589));
    Span4Mux_h I__4568 (
            .O(N__23597),
            .I(N__23584));
    LocalMux I__4567 (
            .O(N__23594),
            .I(N__23584));
    Span4Mux_h I__4566 (
            .O(N__23589),
            .I(N__23581));
    Span4Mux_v I__4565 (
            .O(N__23584),
            .I(N__23578));
    Odrv4 I__4564 (
            .O(N__23581),
            .I(N_1248_0));
    Odrv4 I__4563 (
            .O(N__23578),
            .I(N_1248_0));
    InMux I__4562 (
            .O(N__23573),
            .I(N__23570));
    LocalMux I__4561 (
            .O(N__23570),
            .I(\this_reset_cond.M_stage_qZ0Z_2 ));
    CascadeMux I__4560 (
            .O(N__23567),
            .I(M_this_spr_ram_write_en_0_i_1_0_cascade_));
    CEMux I__4559 (
            .O(N__23564),
            .I(N__23561));
    LocalMux I__4558 (
            .O(N__23561),
            .I(N__23558));
    Span4Mux_h I__4557 (
            .O(N__23558),
            .I(N__23554));
    CEMux I__4556 (
            .O(N__23557),
            .I(N__23551));
    Span4Mux_h I__4555 (
            .O(N__23554),
            .I(N__23548));
    LocalMux I__4554 (
            .O(N__23551),
            .I(N__23545));
    Sp12to4 I__4553 (
            .O(N__23548),
            .I(N__23542));
    Sp12to4 I__4552 (
            .O(N__23545),
            .I(N__23539));
    Span12Mux_v I__4551 (
            .O(N__23542),
            .I(N__23534));
    Span12Mux_v I__4550 (
            .O(N__23539),
            .I(N__23534));
    Odrv12 I__4549 (
            .O(N__23534),
            .I(\this_spr_ram.mem_WE_2 ));
    InMux I__4548 (
            .O(N__23531),
            .I(N__23528));
    LocalMux I__4547 (
            .O(N__23528),
            .I(N__23525));
    Span4Mux_v I__4546 (
            .O(N__23525),
            .I(N__23522));
    Odrv4 I__4545 (
            .O(N__23522),
            .I(\this_vga_signals.M_vcounter_d7lt8_0 ));
    InMux I__4544 (
            .O(N__23519),
            .I(N__23516));
    LocalMux I__4543 (
            .O(N__23516),
            .I(N__23513));
    Span4Mux_h I__4542 (
            .O(N__23513),
            .I(N__23510));
    Span4Mux_h I__4541 (
            .O(N__23510),
            .I(N__23507));
    Span4Mux_h I__4540 (
            .O(N__23507),
            .I(N__23504));
    Odrv4 I__4539 (
            .O(N__23504),
            .I(\this_delay_clk.M_pipe_qZ0Z_3 ));
    CEMux I__4538 (
            .O(N__23501),
            .I(N__23498));
    LocalMux I__4537 (
            .O(N__23498),
            .I(N__23495));
    Span4Mux_h I__4536 (
            .O(N__23495),
            .I(N__23492));
    Odrv4 I__4535 (
            .O(N__23492),
            .I(N_1256_0));
    InMux I__4534 (
            .O(N__23489),
            .I(N__23486));
    LocalMux I__4533 (
            .O(N__23486),
            .I(N__23483));
    Span4Mux_h I__4532 (
            .O(N__23483),
            .I(N__23479));
    InMux I__4531 (
            .O(N__23482),
            .I(N__23476));
    Sp12to4 I__4530 (
            .O(N__23479),
            .I(N__23473));
    LocalMux I__4529 (
            .O(N__23476),
            .I(N__23470));
    Span12Mux_v I__4528 (
            .O(N__23473),
            .I(N__23467));
    Span12Mux_v I__4527 (
            .O(N__23470),
            .I(N__23464));
    Odrv12 I__4526 (
            .O(N__23467),
            .I(M_this_oam_ram_read_data_16));
    Odrv12 I__4525 (
            .O(N__23464),
            .I(M_this_oam_ram_read_data_16));
    InMux I__4524 (
            .O(N__23459),
            .I(N__23456));
    LocalMux I__4523 (
            .O(N__23456),
            .I(N__23453));
    Span4Mux_v I__4522 (
            .O(N__23453),
            .I(N__23450));
    Span4Mux_h I__4521 (
            .O(N__23450),
            .I(N__23447));
    Odrv4 I__4520 (
            .O(N__23447),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_16 ));
    InMux I__4519 (
            .O(N__23444),
            .I(N__23441));
    LocalMux I__4518 (
            .O(N__23441),
            .I(N__23438));
    Span4Mux_v I__4517 (
            .O(N__23438),
            .I(N__23434));
    InMux I__4516 (
            .O(N__23437),
            .I(N__23431));
    Span4Mux_h I__4515 (
            .O(N__23434),
            .I(N__23426));
    LocalMux I__4514 (
            .O(N__23431),
            .I(N__23426));
    Sp12to4 I__4513 (
            .O(N__23426),
            .I(N__23423));
    Span12Mux_v I__4512 (
            .O(N__23423),
            .I(N__23420));
    Odrv12 I__4511 (
            .O(N__23420),
            .I(M_this_oam_ram_read_data_17));
    InMux I__4510 (
            .O(N__23417),
            .I(N__23414));
    LocalMux I__4509 (
            .O(N__23414),
            .I(N__23411));
    Span4Mux_v I__4508 (
            .O(N__23411),
            .I(N__23408));
    Span4Mux_h I__4507 (
            .O(N__23408),
            .I(N__23405));
    Odrv4 I__4506 (
            .O(N__23405),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_17 ));
    InMux I__4505 (
            .O(N__23402),
            .I(N__23399));
    LocalMux I__4504 (
            .O(N__23399),
            .I(N__23395));
    InMux I__4503 (
            .O(N__23398),
            .I(N__23392));
    Span4Mux_h I__4502 (
            .O(N__23395),
            .I(N__23389));
    LocalMux I__4501 (
            .O(N__23392),
            .I(N__23386));
    Sp12to4 I__4500 (
            .O(N__23389),
            .I(N__23383));
    Span4Mux_v I__4499 (
            .O(N__23386),
            .I(N__23380));
    Span12Mux_v I__4498 (
            .O(N__23383),
            .I(N__23377));
    Span4Mux_v I__4497 (
            .O(N__23380),
            .I(N__23374));
    Odrv12 I__4496 (
            .O(N__23377),
            .I(M_this_oam_ram_read_data_18));
    Odrv4 I__4495 (
            .O(N__23374),
            .I(M_this_oam_ram_read_data_18));
    InMux I__4494 (
            .O(N__23369),
            .I(N__23366));
    LocalMux I__4493 (
            .O(N__23366),
            .I(N__23363));
    Span4Mux_h I__4492 (
            .O(N__23363),
            .I(N__23360));
    Span4Mux_h I__4491 (
            .O(N__23360),
            .I(N__23357));
    Odrv4 I__4490 (
            .O(N__23357),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_18 ));
    InMux I__4489 (
            .O(N__23354),
            .I(N__23351));
    LocalMux I__4488 (
            .O(N__23351),
            .I(N__23348));
    Span4Mux_h I__4487 (
            .O(N__23348),
            .I(N__23345));
    Sp12to4 I__4486 (
            .O(N__23345),
            .I(N__23342));
    Span12Mux_v I__4485 (
            .O(N__23342),
            .I(N__23339));
    Odrv12 I__4484 (
            .O(N__23339),
            .I(M_this_oam_ram_read_data_27));
    InMux I__4483 (
            .O(N__23336),
            .I(N__23333));
    LocalMux I__4482 (
            .O(N__23333),
            .I(N__23330));
    Odrv12 I__4481 (
            .O(N__23330),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_27 ));
    InMux I__4480 (
            .O(N__23327),
            .I(\this_ppu.un1_M_surface_y_d_cry_5 ));
    CascadeMux I__4479 (
            .O(N__23324),
            .I(N__23321));
    InMux I__4478 (
            .O(N__23321),
            .I(N__23317));
    CascadeMux I__4477 (
            .O(N__23320),
            .I(N__23314));
    LocalMux I__4476 (
            .O(N__23317),
            .I(N__23311));
    InMux I__4475 (
            .O(N__23314),
            .I(N__23308));
    Odrv12 I__4474 (
            .O(N__23311),
            .I(\this_ppu.M_screen_y_qZ0Z_7 ));
    LocalMux I__4473 (
            .O(N__23308),
            .I(\this_ppu.M_screen_y_qZ0Z_7 ));
    InMux I__4472 (
            .O(N__23303),
            .I(bfn_14_19_0_));
    CascadeMux I__4471 (
            .O(N__23300),
            .I(N__23297));
    CascadeBuf I__4470 (
            .O(N__23297),
            .I(N__23293));
    InMux I__4469 (
            .O(N__23296),
            .I(N__23290));
    CascadeMux I__4468 (
            .O(N__23293),
            .I(N__23287));
    LocalMux I__4467 (
            .O(N__23290),
            .I(N__23284));
    InMux I__4466 (
            .O(N__23287),
            .I(N__23281));
    Span4Mux_v I__4465 (
            .O(N__23284),
            .I(N__23278));
    LocalMux I__4464 (
            .O(N__23281),
            .I(N__23275));
    Span4Mux_h I__4463 (
            .O(N__23278),
            .I(N__23272));
    Span12Mux_h I__4462 (
            .O(N__23275),
            .I(N__23269));
    Odrv4 I__4461 (
            .O(N__23272),
            .I(M_this_ppu_map_addr_9));
    Odrv12 I__4460 (
            .O(N__23269),
            .I(M_this_ppu_map_addr_9));
    CascadeMux I__4459 (
            .O(N__23264),
            .I(N__23261));
    InMux I__4458 (
            .O(N__23261),
            .I(N__23258));
    LocalMux I__4457 (
            .O(N__23258),
            .I(N__23250));
    CascadeMux I__4456 (
            .O(N__23257),
            .I(N__23247));
    InMux I__4455 (
            .O(N__23256),
            .I(N__23242));
    InMux I__4454 (
            .O(N__23255),
            .I(N__23242));
    InMux I__4453 (
            .O(N__23254),
            .I(N__23236));
    InMux I__4452 (
            .O(N__23253),
            .I(N__23236));
    Span12Mux_v I__4451 (
            .O(N__23250),
            .I(N__23233));
    InMux I__4450 (
            .O(N__23247),
            .I(N__23230));
    LocalMux I__4449 (
            .O(N__23242),
            .I(N__23227));
    InMux I__4448 (
            .O(N__23241),
            .I(N__23224));
    LocalMux I__4447 (
            .O(N__23236),
            .I(N__23221));
    Odrv12 I__4446 (
            .O(N__23233),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__4445 (
            .O(N__23230),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__4444 (
            .O(N__23227),
            .I(M_this_ppu_vram_addr_7));
    LocalMux I__4443 (
            .O(N__23224),
            .I(M_this_ppu_vram_addr_7));
    Odrv4 I__4442 (
            .O(N__23221),
            .I(M_this_ppu_vram_addr_7));
    InMux I__4441 (
            .O(N__23210),
            .I(N__23204));
    InMux I__4440 (
            .O(N__23209),
            .I(N__23201));
    InMux I__4439 (
            .O(N__23208),
            .I(N__23196));
    InMux I__4438 (
            .O(N__23207),
            .I(N__23196));
    LocalMux I__4437 (
            .O(N__23204),
            .I(N__23193));
    LocalMux I__4436 (
            .O(N__23201),
            .I(N__23190));
    LocalMux I__4435 (
            .O(N__23196),
            .I(\this_ppu.M_screen_y_qZ0Z_1 ));
    Odrv4 I__4434 (
            .O(N__23193),
            .I(\this_ppu.M_screen_y_qZ0Z_1 ));
    Odrv12 I__4433 (
            .O(N__23190),
            .I(\this_ppu.M_screen_y_qZ0Z_1 ));
    CascadeMux I__4432 (
            .O(N__23183),
            .I(N__23172));
    InMux I__4431 (
            .O(N__23182),
            .I(N__23168));
    InMux I__4430 (
            .O(N__23181),
            .I(N__23159));
    InMux I__4429 (
            .O(N__23180),
            .I(N__23159));
    InMux I__4428 (
            .O(N__23179),
            .I(N__23159));
    InMux I__4427 (
            .O(N__23178),
            .I(N__23159));
    InMux I__4426 (
            .O(N__23177),
            .I(N__23151));
    InMux I__4425 (
            .O(N__23176),
            .I(N__23151));
    InMux I__4424 (
            .O(N__23175),
            .I(N__23151));
    InMux I__4423 (
            .O(N__23172),
            .I(N__23148));
    InMux I__4422 (
            .O(N__23171),
            .I(N__23145));
    LocalMux I__4421 (
            .O(N__23168),
            .I(N__23133));
    LocalMux I__4420 (
            .O(N__23159),
            .I(N__23133));
    InMux I__4419 (
            .O(N__23158),
            .I(N__23130));
    LocalMux I__4418 (
            .O(N__23151),
            .I(N__23123));
    LocalMux I__4417 (
            .O(N__23148),
            .I(N__23123));
    LocalMux I__4416 (
            .O(N__23145),
            .I(N__23123));
    InMux I__4415 (
            .O(N__23144),
            .I(N__23114));
    InMux I__4414 (
            .O(N__23143),
            .I(N__23114));
    InMux I__4413 (
            .O(N__23142),
            .I(N__23114));
    InMux I__4412 (
            .O(N__23141),
            .I(N__23114));
    InMux I__4411 (
            .O(N__23140),
            .I(N__23107));
    InMux I__4410 (
            .O(N__23139),
            .I(N__23107));
    InMux I__4409 (
            .O(N__23138),
            .I(N__23107));
    Odrv4 I__4408 (
            .O(N__23133),
            .I(M_this_ppu_vga_is_drawing));
    LocalMux I__4407 (
            .O(N__23130),
            .I(M_this_ppu_vga_is_drawing));
    Odrv4 I__4406 (
            .O(N__23123),
            .I(M_this_ppu_vga_is_drawing));
    LocalMux I__4405 (
            .O(N__23114),
            .I(M_this_ppu_vga_is_drawing));
    LocalMux I__4404 (
            .O(N__23107),
            .I(M_this_ppu_vga_is_drawing));
    InMux I__4403 (
            .O(N__23096),
            .I(N__23091));
    CascadeMux I__4402 (
            .O(N__23095),
            .I(N__23087));
    InMux I__4401 (
            .O(N__23094),
            .I(N__23084));
    LocalMux I__4400 (
            .O(N__23091),
            .I(N__23081));
    InMux I__4399 (
            .O(N__23090),
            .I(N__23078));
    InMux I__4398 (
            .O(N__23087),
            .I(N__23075));
    LocalMux I__4397 (
            .O(N__23084),
            .I(N__23072));
    Span4Mux_h I__4396 (
            .O(N__23081),
            .I(N__23067));
    LocalMux I__4395 (
            .O(N__23078),
            .I(N__23067));
    LocalMux I__4394 (
            .O(N__23075),
            .I(\this_ppu.M_screen_y_qZ0Z_2 ));
    Odrv12 I__4393 (
            .O(N__23072),
            .I(\this_ppu.M_screen_y_qZ0Z_2 ));
    Odrv4 I__4392 (
            .O(N__23067),
            .I(\this_ppu.M_screen_y_qZ0Z_2 ));
    CEMux I__4391 (
            .O(N__23060),
            .I(N__23055));
    CEMux I__4390 (
            .O(N__23059),
            .I(N__23052));
    CEMux I__4389 (
            .O(N__23058),
            .I(N__23048));
    LocalMux I__4388 (
            .O(N__23055),
            .I(N__23045));
    LocalMux I__4387 (
            .O(N__23052),
            .I(N__23042));
    CEMux I__4386 (
            .O(N__23051),
            .I(N__23039));
    LocalMux I__4385 (
            .O(N__23048),
            .I(N__23036));
    Span4Mux_v I__4384 (
            .O(N__23045),
            .I(N__23029));
    Span4Mux_v I__4383 (
            .O(N__23042),
            .I(N__23029));
    LocalMux I__4382 (
            .O(N__23039),
            .I(N__23029));
    Span4Mux_h I__4381 (
            .O(N__23036),
            .I(N__23026));
    Odrv4 I__4380 (
            .O(N__23029),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0 ));
    Odrv4 I__4379 (
            .O(N__23026),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0 ));
    InMux I__4378 (
            .O(N__23021),
            .I(N__23018));
    LocalMux I__4377 (
            .O(N__23018),
            .I(N__23015));
    Span12Mux_h I__4376 (
            .O(N__23015),
            .I(N__23012));
    Odrv12 I__4375 (
            .O(N__23012),
            .I(M_this_oam_ram_read_data_12));
    InMux I__4374 (
            .O(N__23009),
            .I(N__23006));
    LocalMux I__4373 (
            .O(N__23006),
            .I(N__23003));
    Span4Mux_h I__4372 (
            .O(N__23003),
            .I(N__23000));
    Span4Mux_h I__4371 (
            .O(N__23000),
            .I(N__22997));
    Odrv4 I__4370 (
            .O(N__22997),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_12 ));
    CascadeMux I__4369 (
            .O(N__22994),
            .I(N__22990));
    CascadeMux I__4368 (
            .O(N__22993),
            .I(N__22984));
    InMux I__4367 (
            .O(N__22990),
            .I(N__22979));
    CascadeMux I__4366 (
            .O(N__22989),
            .I(N__22976));
    CascadeMux I__4365 (
            .O(N__22988),
            .I(N__22973));
    CascadeMux I__4364 (
            .O(N__22987),
            .I(N__22968));
    InMux I__4363 (
            .O(N__22984),
            .I(N__22964));
    CascadeMux I__4362 (
            .O(N__22983),
            .I(N__22961));
    CascadeMux I__4361 (
            .O(N__22982),
            .I(N__22958));
    LocalMux I__4360 (
            .O(N__22979),
            .I(N__22954));
    InMux I__4359 (
            .O(N__22976),
            .I(N__22951));
    InMux I__4358 (
            .O(N__22973),
            .I(N__22948));
    CascadeMux I__4357 (
            .O(N__22972),
            .I(N__22945));
    CascadeMux I__4356 (
            .O(N__22971),
            .I(N__22942));
    InMux I__4355 (
            .O(N__22968),
            .I(N__22937));
    CascadeMux I__4354 (
            .O(N__22967),
            .I(N__22934));
    LocalMux I__4353 (
            .O(N__22964),
            .I(N__22931));
    InMux I__4352 (
            .O(N__22961),
            .I(N__22928));
    InMux I__4351 (
            .O(N__22958),
            .I(N__22925));
    CascadeMux I__4350 (
            .O(N__22957),
            .I(N__22922));
    Span4Mux_s0_v I__4349 (
            .O(N__22954),
            .I(N__22916));
    LocalMux I__4348 (
            .O(N__22951),
            .I(N__22916));
    LocalMux I__4347 (
            .O(N__22948),
            .I(N__22913));
    InMux I__4346 (
            .O(N__22945),
            .I(N__22910));
    InMux I__4345 (
            .O(N__22942),
            .I(N__22907));
    CascadeMux I__4344 (
            .O(N__22941),
            .I(N__22904));
    CascadeMux I__4343 (
            .O(N__22940),
            .I(N__22901));
    LocalMux I__4342 (
            .O(N__22937),
            .I(N__22897));
    InMux I__4341 (
            .O(N__22934),
            .I(N__22894));
    Span4Mux_h I__4340 (
            .O(N__22931),
            .I(N__22891));
    LocalMux I__4339 (
            .O(N__22928),
            .I(N__22888));
    LocalMux I__4338 (
            .O(N__22925),
            .I(N__22885));
    InMux I__4337 (
            .O(N__22922),
            .I(N__22882));
    CascadeMux I__4336 (
            .O(N__22921),
            .I(N__22879));
    Span4Mux_v I__4335 (
            .O(N__22916),
            .I(N__22872));
    Span4Mux_h I__4334 (
            .O(N__22913),
            .I(N__22872));
    LocalMux I__4333 (
            .O(N__22910),
            .I(N__22872));
    LocalMux I__4332 (
            .O(N__22907),
            .I(N__22869));
    InMux I__4331 (
            .O(N__22904),
            .I(N__22866));
    InMux I__4330 (
            .O(N__22901),
            .I(N__22863));
    CascadeMux I__4329 (
            .O(N__22900),
            .I(N__22860));
    Span4Mux_h I__4328 (
            .O(N__22897),
            .I(N__22856));
    LocalMux I__4327 (
            .O(N__22894),
            .I(N__22853));
    Span4Mux_v I__4326 (
            .O(N__22891),
            .I(N__22848));
    Span4Mux_h I__4325 (
            .O(N__22888),
            .I(N__22848));
    Span4Mux_h I__4324 (
            .O(N__22885),
            .I(N__22845));
    LocalMux I__4323 (
            .O(N__22882),
            .I(N__22842));
    InMux I__4322 (
            .O(N__22879),
            .I(N__22839));
    Span4Mux_v I__4321 (
            .O(N__22872),
            .I(N__22832));
    Span4Mux_h I__4320 (
            .O(N__22869),
            .I(N__22832));
    LocalMux I__4319 (
            .O(N__22866),
            .I(N__22832));
    LocalMux I__4318 (
            .O(N__22863),
            .I(N__22829));
    InMux I__4317 (
            .O(N__22860),
            .I(N__22826));
    CascadeMux I__4316 (
            .O(N__22859),
            .I(N__22823));
    Span4Mux_h I__4315 (
            .O(N__22856),
            .I(N__22820));
    Span4Mux_h I__4314 (
            .O(N__22853),
            .I(N__22817));
    Span4Mux_v I__4313 (
            .O(N__22848),
            .I(N__22814));
    Span4Mux_v I__4312 (
            .O(N__22845),
            .I(N__22809));
    Span4Mux_h I__4311 (
            .O(N__22842),
            .I(N__22809));
    LocalMux I__4310 (
            .O(N__22839),
            .I(N__22806));
    Span4Mux_v I__4309 (
            .O(N__22832),
            .I(N__22799));
    Span4Mux_h I__4308 (
            .O(N__22829),
            .I(N__22799));
    LocalMux I__4307 (
            .O(N__22826),
            .I(N__22799));
    InMux I__4306 (
            .O(N__22823),
            .I(N__22796));
    Sp12to4 I__4305 (
            .O(N__22820),
            .I(N__22793));
    Span4Mux_h I__4304 (
            .O(N__22817),
            .I(N__22790));
    Span4Mux_v I__4303 (
            .O(N__22814),
            .I(N__22787));
    Span4Mux_h I__4302 (
            .O(N__22809),
            .I(N__22784));
    Span12Mux_s10_h I__4301 (
            .O(N__22806),
            .I(N__22781));
    Span4Mux_v I__4300 (
            .O(N__22799),
            .I(N__22778));
    LocalMux I__4299 (
            .O(N__22796),
            .I(N__22775));
    Span12Mux_s11_v I__4298 (
            .O(N__22793),
            .I(N__22770));
    Sp12to4 I__4297 (
            .O(N__22790),
            .I(N__22770));
    Span4Mux_h I__4296 (
            .O(N__22787),
            .I(N__22765));
    Span4Mux_v I__4295 (
            .O(N__22784),
            .I(N__22765));
    Span12Mux_v I__4294 (
            .O(N__22781),
            .I(N__22758));
    Sp12to4 I__4293 (
            .O(N__22778),
            .I(N__22758));
    Span12Mux_s9_h I__4292 (
            .O(N__22775),
            .I(N__22758));
    Odrv12 I__4291 (
            .O(N__22770),
            .I(M_this_ppu_spr_addr_8));
    Odrv4 I__4290 (
            .O(N__22765),
            .I(M_this_ppu_spr_addr_8));
    Odrv12 I__4289 (
            .O(N__22758),
            .I(M_this_ppu_spr_addr_8));
    InMux I__4288 (
            .O(N__22751),
            .I(N__22748));
    LocalMux I__4287 (
            .O(N__22748),
            .I(N__22745));
    Odrv4 I__4286 (
            .O(N__22745),
            .I(\this_ppu.M_screen_y_q_RNICCMV8Z0Z_0 ));
    CascadeMux I__4285 (
            .O(N__22742),
            .I(N__22738));
    InMux I__4284 (
            .O(N__22741),
            .I(N__22734));
    InMux I__4283 (
            .O(N__22738),
            .I(N__22731));
    InMux I__4282 (
            .O(N__22737),
            .I(N__22728));
    LocalMux I__4281 (
            .O(N__22734),
            .I(N__22723));
    LocalMux I__4280 (
            .O(N__22731),
            .I(N__22723));
    LocalMux I__4279 (
            .O(N__22728),
            .I(N__22720));
    Span4Mux_v I__4278 (
            .O(N__22723),
            .I(N__22717));
    Span4Mux_v I__4277 (
            .O(N__22720),
            .I(N__22714));
    Span4Mux_h I__4276 (
            .O(N__22717),
            .I(N__22711));
    Odrv4 I__4275 (
            .O(N__22714),
            .I(\this_ppu.offset_y ));
    Odrv4 I__4274 (
            .O(N__22711),
            .I(\this_ppu.offset_y ));
    InMux I__4273 (
            .O(N__22706),
            .I(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ));
    InMux I__4272 (
            .O(N__22703),
            .I(N__22700));
    LocalMux I__4271 (
            .O(N__22700),
            .I(N__22697));
    Odrv4 I__4270 (
            .O(N__22697),
            .I(\this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1 ));
    CascadeMux I__4269 (
            .O(N__22694),
            .I(N__22690));
    InMux I__4268 (
            .O(N__22693),
            .I(N__22687));
    InMux I__4267 (
            .O(N__22690),
            .I(N__22684));
    LocalMux I__4266 (
            .O(N__22687),
            .I(N__22681));
    LocalMux I__4265 (
            .O(N__22684),
            .I(N__22678));
    Span4Mux_v I__4264 (
            .O(N__22681),
            .I(N__22673));
    Span4Mux_h I__4263 (
            .O(N__22678),
            .I(N__22673));
    Span4Mux_h I__4262 (
            .O(N__22673),
            .I(N__22670));
    Odrv4 I__4261 (
            .O(N__22670),
            .I(\this_ppu.M_surface_y_qZ0Z_1 ));
    InMux I__4260 (
            .O(N__22667),
            .I(\this_ppu.un1_M_surface_y_d_cry_0 ));
    InMux I__4259 (
            .O(N__22664),
            .I(N__22661));
    LocalMux I__4258 (
            .O(N__22661),
            .I(N__22658));
    Span4Mux_v I__4257 (
            .O(N__22658),
            .I(N__22655));
    Odrv4 I__4256 (
            .O(N__22655),
            .I(\this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2 ));
    CascadeMux I__4255 (
            .O(N__22652),
            .I(N__22648));
    InMux I__4254 (
            .O(N__22651),
            .I(N__22645));
    InMux I__4253 (
            .O(N__22648),
            .I(N__22642));
    LocalMux I__4252 (
            .O(N__22645),
            .I(N__22639));
    LocalMux I__4251 (
            .O(N__22642),
            .I(N__22636));
    Span4Mux_h I__4250 (
            .O(N__22639),
            .I(N__22633));
    Span12Mux_h I__4249 (
            .O(N__22636),
            .I(N__22630));
    Odrv4 I__4248 (
            .O(N__22633),
            .I(\this_ppu.M_surface_y_qZ0Z_2 ));
    Odrv12 I__4247 (
            .O(N__22630),
            .I(\this_ppu.M_surface_y_qZ0Z_2 ));
    InMux I__4246 (
            .O(N__22625),
            .I(\this_ppu.un1_M_surface_y_d_cry_1 ));
    InMux I__4245 (
            .O(N__22622),
            .I(N__22619));
    LocalMux I__4244 (
            .O(N__22619),
            .I(N__22616));
    Odrv4 I__4243 (
            .O(N__22616),
            .I(\this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3 ));
    CascadeMux I__4242 (
            .O(N__22613),
            .I(N__22610));
    CascadeBuf I__4241 (
            .O(N__22610),
            .I(N__22607));
    CascadeMux I__4240 (
            .O(N__22607),
            .I(N__22603));
    CascadeMux I__4239 (
            .O(N__22606),
            .I(N__22600));
    InMux I__4238 (
            .O(N__22603),
            .I(N__22597));
    InMux I__4237 (
            .O(N__22600),
            .I(N__22594));
    LocalMux I__4236 (
            .O(N__22597),
            .I(N__22591));
    LocalMux I__4235 (
            .O(N__22594),
            .I(N__22588));
    Span4Mux_v I__4234 (
            .O(N__22591),
            .I(N__22585));
    Span4Mux_h I__4233 (
            .O(N__22588),
            .I(N__22582));
    Sp12to4 I__4232 (
            .O(N__22585),
            .I(N__22579));
    Span4Mux_h I__4231 (
            .O(N__22582),
            .I(N__22576));
    Span12Mux_v I__4230 (
            .O(N__22579),
            .I(N__22573));
    Odrv4 I__4229 (
            .O(N__22576),
            .I(M_this_ppu_map_addr_5));
    Odrv12 I__4228 (
            .O(N__22573),
            .I(M_this_ppu_map_addr_5));
    InMux I__4227 (
            .O(N__22568),
            .I(\this_ppu.un1_M_surface_y_d_cry_2 ));
    InMux I__4226 (
            .O(N__22565),
            .I(N__22562));
    LocalMux I__4225 (
            .O(N__22562),
            .I(N__22559));
    Odrv4 I__4224 (
            .O(N__22559),
            .I(\this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4 ));
    CascadeMux I__4223 (
            .O(N__22556),
            .I(N__22552));
    CascadeMux I__4222 (
            .O(N__22555),
            .I(N__22549));
    CascadeBuf I__4221 (
            .O(N__22552),
            .I(N__22546));
    InMux I__4220 (
            .O(N__22549),
            .I(N__22543));
    CascadeMux I__4219 (
            .O(N__22546),
            .I(N__22540));
    LocalMux I__4218 (
            .O(N__22543),
            .I(N__22537));
    InMux I__4217 (
            .O(N__22540),
            .I(N__22534));
    Span4Mux_h I__4216 (
            .O(N__22537),
            .I(N__22531));
    LocalMux I__4215 (
            .O(N__22534),
            .I(N__22528));
    Span4Mux_h I__4214 (
            .O(N__22531),
            .I(N__22525));
    Span12Mux_v I__4213 (
            .O(N__22528),
            .I(N__22522));
    Odrv4 I__4212 (
            .O(N__22525),
            .I(M_this_ppu_map_addr_6));
    Odrv12 I__4211 (
            .O(N__22522),
            .I(M_this_ppu_map_addr_6));
    InMux I__4210 (
            .O(N__22517),
            .I(\this_ppu.un1_M_surface_y_d_cry_3 ));
    InMux I__4209 (
            .O(N__22514),
            .I(N__22511));
    LocalMux I__4208 (
            .O(N__22511),
            .I(N__22508));
    Odrv4 I__4207 (
            .O(N__22508),
            .I(\this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5 ));
    CascadeMux I__4206 (
            .O(N__22505),
            .I(N__22502));
    CascadeBuf I__4205 (
            .O(N__22502),
            .I(N__22499));
    CascadeMux I__4204 (
            .O(N__22499),
            .I(N__22496));
    InMux I__4203 (
            .O(N__22496),
            .I(N__22492));
    CascadeMux I__4202 (
            .O(N__22495),
            .I(N__22489));
    LocalMux I__4201 (
            .O(N__22492),
            .I(N__22486));
    InMux I__4200 (
            .O(N__22489),
            .I(N__22483));
    Span4Mux_v I__4199 (
            .O(N__22486),
            .I(N__22480));
    LocalMux I__4198 (
            .O(N__22483),
            .I(N__22477));
    Span4Mux_v I__4197 (
            .O(N__22480),
            .I(N__22474));
    Span4Mux_h I__4196 (
            .O(N__22477),
            .I(N__22471));
    Span4Mux_v I__4195 (
            .O(N__22474),
            .I(N__22468));
    Span4Mux_h I__4194 (
            .O(N__22471),
            .I(N__22465));
    Sp12to4 I__4193 (
            .O(N__22468),
            .I(N__22462));
    Odrv4 I__4192 (
            .O(N__22465),
            .I(M_this_ppu_map_addr_7));
    Odrv12 I__4191 (
            .O(N__22462),
            .I(M_this_ppu_map_addr_7));
    InMux I__4190 (
            .O(N__22457),
            .I(\this_ppu.un1_M_surface_y_d_cry_4 ));
    InMux I__4189 (
            .O(N__22454),
            .I(N__22451));
    LocalMux I__4188 (
            .O(N__22451),
            .I(N__22448));
    Odrv4 I__4187 (
            .O(N__22448),
            .I(\this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6 ));
    CascadeMux I__4186 (
            .O(N__22445),
            .I(N__22442));
    CascadeBuf I__4185 (
            .O(N__22442),
            .I(N__22439));
    CascadeMux I__4184 (
            .O(N__22439),
            .I(N__22435));
    CascadeMux I__4183 (
            .O(N__22438),
            .I(N__22432));
    InMux I__4182 (
            .O(N__22435),
            .I(N__22429));
    InMux I__4181 (
            .O(N__22432),
            .I(N__22426));
    LocalMux I__4180 (
            .O(N__22429),
            .I(N__22423));
    LocalMux I__4179 (
            .O(N__22426),
            .I(N__22420));
    Sp12to4 I__4178 (
            .O(N__22423),
            .I(N__22417));
    Span4Mux_h I__4177 (
            .O(N__22420),
            .I(N__22414));
    Span12Mux_s7_v I__4176 (
            .O(N__22417),
            .I(N__22411));
    Span4Mux_h I__4175 (
            .O(N__22414),
            .I(N__22408));
    Span12Mux_h I__4174 (
            .O(N__22411),
            .I(N__22405));
    Odrv4 I__4173 (
            .O(N__22408),
            .I(M_this_ppu_map_addr_8));
    Odrv12 I__4172 (
            .O(N__22405),
            .I(M_this_ppu_map_addr_8));
    CascadeMux I__4171 (
            .O(N__22400),
            .I(M_this_ppu_vga_is_drawing_cascade_));
    InMux I__4170 (
            .O(N__22397),
            .I(N__22393));
    CascadeMux I__4169 (
            .O(N__22396),
            .I(N__22389));
    LocalMux I__4168 (
            .O(N__22393),
            .I(N__22386));
    InMux I__4167 (
            .O(N__22392),
            .I(N__22382));
    InMux I__4166 (
            .O(N__22389),
            .I(N__22379));
    Span4Mux_h I__4165 (
            .O(N__22386),
            .I(N__22376));
    InMux I__4164 (
            .O(N__22385),
            .I(N__22373));
    LocalMux I__4163 (
            .O(N__22382),
            .I(N__22370));
    LocalMux I__4162 (
            .O(N__22379),
            .I(this_ppu_M_screen_y_q_5));
    Odrv4 I__4161 (
            .O(N__22376),
            .I(this_ppu_M_screen_y_q_5));
    LocalMux I__4160 (
            .O(N__22373),
            .I(this_ppu_M_screen_y_q_5));
    Odrv4 I__4159 (
            .O(N__22370),
            .I(this_ppu_M_screen_y_q_5));
    InMux I__4158 (
            .O(N__22361),
            .I(N__22358));
    LocalMux I__4157 (
            .O(N__22358),
            .I(N__22352));
    InMux I__4156 (
            .O(N__22357),
            .I(N__22349));
    InMux I__4155 (
            .O(N__22356),
            .I(N__22344));
    InMux I__4154 (
            .O(N__22355),
            .I(N__22344));
    Span4Mux_h I__4153 (
            .O(N__22352),
            .I(N__22339));
    LocalMux I__4152 (
            .O(N__22349),
            .I(N__22339));
    LocalMux I__4151 (
            .O(N__22344),
            .I(this_ppu_M_screen_y_q_6));
    Odrv4 I__4150 (
            .O(N__22339),
            .I(this_ppu_M_screen_y_q_6));
    InMux I__4149 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__4148 (
            .O(N__22331),
            .I(\this_ppu.un1_M_surface_x_q_c1 ));
    CascadeMux I__4147 (
            .O(N__22328),
            .I(N__22325));
    InMux I__4146 (
            .O(N__22325),
            .I(N__22322));
    LocalMux I__4145 (
            .O(N__22322),
            .I(N__22319));
    Span4Mux_v I__4144 (
            .O(N__22319),
            .I(N__22316));
    Odrv4 I__4143 (
            .O(N__22316),
            .I(M_this_scroll_qZ0Z_9));
    CascadeMux I__4142 (
            .O(N__22313),
            .I(N__22310));
    InMux I__4141 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__4140 (
            .O(N__22307),
            .I(M_this_scroll_qZ0Z_15));
    InMux I__4139 (
            .O(N__22304),
            .I(N__22301));
    LocalMux I__4138 (
            .O(N__22301),
            .I(N__22298));
    Odrv4 I__4137 (
            .O(N__22298),
            .I(\this_ppu.un1_M_surface_x_q_ac0_11 ));
    InMux I__4136 (
            .O(N__22295),
            .I(N__22292));
    LocalMux I__4135 (
            .O(N__22292),
            .I(N__22289));
    Odrv4 I__4134 (
            .O(N__22289),
            .I(M_this_scroll_qZ0Z_12));
    InMux I__4133 (
            .O(N__22286),
            .I(N__22282));
    InMux I__4132 (
            .O(N__22285),
            .I(N__22279));
    LocalMux I__4131 (
            .O(N__22282),
            .I(\this_ppu.un1_M_surface_x_q_c4 ));
    LocalMux I__4130 (
            .O(N__22279),
            .I(\this_ppu.un1_M_surface_x_q_c4 ));
    CascadeMux I__4129 (
            .O(N__22274),
            .I(N__22271));
    InMux I__4128 (
            .O(N__22271),
            .I(N__22263));
    InMux I__4127 (
            .O(N__22270),
            .I(N__22258));
    InMux I__4126 (
            .O(N__22269),
            .I(N__22258));
    InMux I__4125 (
            .O(N__22268),
            .I(N__22244));
    InMux I__4124 (
            .O(N__22267),
            .I(N__22244));
    InMux I__4123 (
            .O(N__22266),
            .I(N__22241));
    LocalMux I__4122 (
            .O(N__22263),
            .I(N__22236));
    LocalMux I__4121 (
            .O(N__22258),
            .I(N__22236));
    InMux I__4120 (
            .O(N__22257),
            .I(N__22225));
    InMux I__4119 (
            .O(N__22256),
            .I(N__22225));
    InMux I__4118 (
            .O(N__22255),
            .I(N__22225));
    InMux I__4117 (
            .O(N__22254),
            .I(N__22225));
    InMux I__4116 (
            .O(N__22253),
            .I(N__22225));
    InMux I__4115 (
            .O(N__22252),
            .I(N__22220));
    InMux I__4114 (
            .O(N__22251),
            .I(N__22220));
    InMux I__4113 (
            .O(N__22250),
            .I(N__22215));
    InMux I__4112 (
            .O(N__22249),
            .I(N__22215));
    LocalMux I__4111 (
            .O(N__22244),
            .I(N__22210));
    LocalMux I__4110 (
            .O(N__22241),
            .I(N__22210));
    Span4Mux_v I__4109 (
            .O(N__22236),
            .I(N__22207));
    LocalMux I__4108 (
            .O(N__22225),
            .I(N__22204));
    LocalMux I__4107 (
            .O(N__22220),
            .I(N__22199));
    LocalMux I__4106 (
            .O(N__22215),
            .I(N__22199));
    Odrv4 I__4105 (
            .O(N__22210),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ));
    Odrv4 I__4104 (
            .O(N__22207),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ));
    Odrv4 I__4103 (
            .O(N__22204),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ));
    Odrv4 I__4102 (
            .O(N__22199),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ));
    InMux I__4101 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__4100 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_h I__4099 (
            .O(N__22184),
            .I(N__22181));
    Odrv4 I__4098 (
            .O(N__22181),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_2 ));
    InMux I__4097 (
            .O(N__22178),
            .I(N__22175));
    LocalMux I__4096 (
            .O(N__22175),
            .I(N__22172));
    Sp12to4 I__4095 (
            .O(N__22172),
            .I(N__22169));
    Span12Mux_v I__4094 (
            .O(N__22169),
            .I(N__22166));
    Odrv12 I__4093 (
            .O(N__22166),
            .I(M_this_map_ram_read_data_2));
    InMux I__4092 (
            .O(N__22163),
            .I(N__22159));
    InMux I__4091 (
            .O(N__22162),
            .I(N__22156));
    LocalMux I__4090 (
            .O(N__22159),
            .I(\this_ppu.un3_M_screen_y_d_0_c6 ));
    LocalMux I__4089 (
            .O(N__22156),
            .I(\this_ppu.un3_M_screen_y_d_0_c6 ));
    InMux I__4088 (
            .O(N__22151),
            .I(N__22147));
    InMux I__4087 (
            .O(N__22150),
            .I(N__22144));
    LocalMux I__4086 (
            .O(N__22147),
            .I(N__22141));
    LocalMux I__4085 (
            .O(N__22144),
            .I(\this_ppu.un3_M_screen_y_d_0_c4 ));
    Odrv4 I__4084 (
            .O(N__22141),
            .I(\this_ppu.un3_M_screen_y_d_0_c4 ));
    InMux I__4083 (
            .O(N__22136),
            .I(N__22131));
    InMux I__4082 (
            .O(N__22135),
            .I(N__22128));
    CascadeMux I__4081 (
            .O(N__22134),
            .I(N__22125));
    LocalMux I__4080 (
            .O(N__22131),
            .I(N__22120));
    LocalMux I__4079 (
            .O(N__22128),
            .I(N__22120));
    InMux I__4078 (
            .O(N__22125),
            .I(N__22115));
    Span4Mux_v I__4077 (
            .O(N__22120),
            .I(N__22112));
    InMux I__4076 (
            .O(N__22119),
            .I(N__22109));
    InMux I__4075 (
            .O(N__22118),
            .I(N__22106));
    LocalMux I__4074 (
            .O(N__22115),
            .I(this_ppu_M_screen_y_q_3));
    Odrv4 I__4073 (
            .O(N__22112),
            .I(this_ppu_M_screen_y_q_3));
    LocalMux I__4072 (
            .O(N__22109),
            .I(this_ppu_M_screen_y_q_3));
    LocalMux I__4071 (
            .O(N__22106),
            .I(this_ppu_M_screen_y_q_3));
    InMux I__4070 (
            .O(N__22097),
            .I(N__22093));
    InMux I__4069 (
            .O(N__22096),
            .I(N__22090));
    LocalMux I__4068 (
            .O(N__22093),
            .I(\this_ppu.un3_M_screen_y_d_0_c2 ));
    LocalMux I__4067 (
            .O(N__22090),
            .I(\this_ppu.un3_M_screen_y_d_0_c2 ));
    InMux I__4066 (
            .O(N__22085),
            .I(N__22081));
    InMux I__4065 (
            .O(N__22084),
            .I(N__22078));
    LocalMux I__4064 (
            .O(N__22081),
            .I(N__22072));
    LocalMux I__4063 (
            .O(N__22078),
            .I(N__22069));
    InMux I__4062 (
            .O(N__22077),
            .I(N__22066));
    InMux I__4061 (
            .O(N__22076),
            .I(N__22063));
    InMux I__4060 (
            .O(N__22075),
            .I(N__22060));
    Span4Mux_h I__4059 (
            .O(N__22072),
            .I(N__22057));
    Span4Mux_v I__4058 (
            .O(N__22069),
            .I(N__22054));
    LocalMux I__4057 (
            .O(N__22066),
            .I(this_ppu_M_screen_y_q_4));
    LocalMux I__4056 (
            .O(N__22063),
            .I(this_ppu_M_screen_y_q_4));
    LocalMux I__4055 (
            .O(N__22060),
            .I(this_ppu_M_screen_y_q_4));
    Odrv4 I__4054 (
            .O(N__22057),
            .I(this_ppu_M_screen_y_q_4));
    Odrv4 I__4053 (
            .O(N__22054),
            .I(this_ppu_M_screen_y_q_4));
    InMux I__4052 (
            .O(N__22043),
            .I(N__22038));
    InMux I__4051 (
            .O(N__22042),
            .I(N__22035));
    InMux I__4050 (
            .O(N__22041),
            .I(N__22032));
    LocalMux I__4049 (
            .O(N__22038),
            .I(N__22029));
    LocalMux I__4048 (
            .O(N__22035),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    LocalMux I__4047 (
            .O(N__22032),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    Odrv4 I__4046 (
            .O(N__22029),
            .I(\this_ppu.M_state_qZ0Z_6 ));
    CascadeMux I__4045 (
            .O(N__22022),
            .I(\this_ppu.m68_0_a2_2_cascade_ ));
    InMux I__4044 (
            .O(N__22019),
            .I(N__22016));
    LocalMux I__4043 (
            .O(N__22016),
            .I(N__22012));
    InMux I__4042 (
            .O(N__22015),
            .I(N__22009));
    Span4Mux_h I__4041 (
            .O(N__22012),
            .I(N__22006));
    LocalMux I__4040 (
            .O(N__22009),
            .I(N__22003));
    Odrv4 I__4039 (
            .O(N__22006),
            .I(\this_ppu.M_state_q_ns_7 ));
    Odrv4 I__4038 (
            .O(N__22003),
            .I(\this_ppu.M_state_q_ns_7 ));
    CascadeMux I__4037 (
            .O(N__21998),
            .I(N__21995));
    InMux I__4036 (
            .O(N__21995),
            .I(N__21986));
    InMux I__4035 (
            .O(N__21994),
            .I(N__21986));
    InMux I__4034 (
            .O(N__21993),
            .I(N__21981));
    InMux I__4033 (
            .O(N__21992),
            .I(N__21981));
    InMux I__4032 (
            .O(N__21991),
            .I(N__21973));
    LocalMux I__4031 (
            .O(N__21986),
            .I(N__21968));
    LocalMux I__4030 (
            .O(N__21981),
            .I(N__21968));
    InMux I__4029 (
            .O(N__21980),
            .I(N__21957));
    InMux I__4028 (
            .O(N__21979),
            .I(N__21957));
    InMux I__4027 (
            .O(N__21978),
            .I(N__21957));
    InMux I__4026 (
            .O(N__21977),
            .I(N__21957));
    InMux I__4025 (
            .O(N__21976),
            .I(N__21957));
    LocalMux I__4024 (
            .O(N__21973),
            .I(\this_ppu.N_814 ));
    Odrv4 I__4023 (
            .O(N__21968),
            .I(\this_ppu.N_814 ));
    LocalMux I__4022 (
            .O(N__21957),
            .I(\this_ppu.N_814 ));
    InMux I__4021 (
            .O(N__21950),
            .I(N__21939));
    InMux I__4020 (
            .O(N__21949),
            .I(N__21936));
    InMux I__4019 (
            .O(N__21948),
            .I(N__21931));
    InMux I__4018 (
            .O(N__21947),
            .I(N__21931));
    InMux I__4017 (
            .O(N__21946),
            .I(N__21928));
    InMux I__4016 (
            .O(N__21945),
            .I(N__21919));
    InMux I__4015 (
            .O(N__21944),
            .I(N__21919));
    InMux I__4014 (
            .O(N__21943),
            .I(N__21919));
    InMux I__4013 (
            .O(N__21942),
            .I(N__21919));
    LocalMux I__4012 (
            .O(N__21939),
            .I(\this_ppu.N_783 ));
    LocalMux I__4011 (
            .O(N__21936),
            .I(\this_ppu.N_783 ));
    LocalMux I__4010 (
            .O(N__21931),
            .I(\this_ppu.N_783 ));
    LocalMux I__4009 (
            .O(N__21928),
            .I(\this_ppu.N_783 ));
    LocalMux I__4008 (
            .O(N__21919),
            .I(\this_ppu.N_783 ));
    CascadeMux I__4007 (
            .O(N__21908),
            .I(N__21905));
    InMux I__4006 (
            .O(N__21905),
            .I(N__21902));
    LocalMux I__4005 (
            .O(N__21902),
            .I(\this_ppu.M_state_q_RNISP3R6_3Z0Z_10 ));
    InMux I__4004 (
            .O(N__21899),
            .I(N__21894));
    InMux I__4003 (
            .O(N__21898),
            .I(N__21889));
    InMux I__4002 (
            .O(N__21897),
            .I(N__21889));
    LocalMux I__4001 (
            .O(N__21894),
            .I(N__21886));
    LocalMux I__4000 (
            .O(N__21889),
            .I(un1_M_this_oam_address_q_c2));
    Odrv4 I__3999 (
            .O(N__21886),
            .I(un1_M_this_oam_address_q_c2));
    InMux I__3998 (
            .O(N__21881),
            .I(N__21878));
    LocalMux I__3997 (
            .O(N__21878),
            .I(N__21875));
    Span4Mux_h I__3996 (
            .O(N__21875),
            .I(N__21872));
    Odrv4 I__3995 (
            .O(N__21872),
            .I(M_this_data_tmp_qZ0Z_18));
    InMux I__3994 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__3993 (
            .O(N__21866),
            .I(N__21863));
    Odrv4 I__3992 (
            .O(N__21863),
            .I(M_this_data_tmp_qZ0Z_1));
    InMux I__3991 (
            .O(N__21860),
            .I(N__21857));
    LocalMux I__3990 (
            .O(N__21857),
            .I(N__21854));
    Odrv4 I__3989 (
            .O(N__21854),
            .I(M_this_data_tmp_qZ0Z_19));
    CEMux I__3988 (
            .O(N__21851),
            .I(N__21845));
    CEMux I__3987 (
            .O(N__21850),
            .I(N__21842));
    CEMux I__3986 (
            .O(N__21849),
            .I(N__21839));
    CEMux I__3985 (
            .O(N__21848),
            .I(N__21836));
    LocalMux I__3984 (
            .O(N__21845),
            .I(N__21831));
    LocalMux I__3983 (
            .O(N__21842),
            .I(N__21831));
    LocalMux I__3982 (
            .O(N__21839),
            .I(N__21826));
    LocalMux I__3981 (
            .O(N__21836),
            .I(N__21826));
    Span4Mux_v I__3980 (
            .O(N__21831),
            .I(N__21821));
    Span4Mux_v I__3979 (
            .O(N__21826),
            .I(N__21818));
    CEMux I__3978 (
            .O(N__21825),
            .I(N__21815));
    CEMux I__3977 (
            .O(N__21824),
            .I(N__21812));
    Odrv4 I__3976 (
            .O(N__21821),
            .I(N_1232_0));
    Odrv4 I__3975 (
            .O(N__21818),
            .I(N_1232_0));
    LocalMux I__3974 (
            .O(N__21815),
            .I(N_1232_0));
    LocalMux I__3973 (
            .O(N__21812),
            .I(N_1232_0));
    InMux I__3972 (
            .O(N__21803),
            .I(N__21800));
    LocalMux I__3971 (
            .O(N__21800),
            .I(\this_ppu.M_state_q_RNISP3R6_2Z0Z_10 ));
    InMux I__3970 (
            .O(N__21797),
            .I(N__21794));
    LocalMux I__3969 (
            .O(N__21794),
            .I(\this_ppu.M_state_q_RNISP3R6_4Z0Z_10 ));
    InMux I__3968 (
            .O(N__21791),
            .I(N__21788));
    LocalMux I__3967 (
            .O(N__21788),
            .I(\this_ppu.M_state_q_RNISP3R6_0Z0Z_10 ));
    InMux I__3966 (
            .O(N__21785),
            .I(N__21781));
    InMux I__3965 (
            .O(N__21784),
            .I(N__21773));
    LocalMux I__3964 (
            .O(N__21781),
            .I(N__21769));
    InMux I__3963 (
            .O(N__21780),
            .I(N__21766));
    InMux I__3962 (
            .O(N__21779),
            .I(N__21763));
    CascadeMux I__3961 (
            .O(N__21778),
            .I(N__21760));
    InMux I__3960 (
            .O(N__21777),
            .I(N__21755));
    InMux I__3959 (
            .O(N__21776),
            .I(N__21755));
    LocalMux I__3958 (
            .O(N__21773),
            .I(N__21752));
    InMux I__3957 (
            .O(N__21772),
            .I(N__21749));
    Span4Mux_v I__3956 (
            .O(N__21769),
            .I(N__21744));
    LocalMux I__3955 (
            .O(N__21766),
            .I(N__21744));
    LocalMux I__3954 (
            .O(N__21763),
            .I(N__21741));
    InMux I__3953 (
            .O(N__21760),
            .I(N__21738));
    LocalMux I__3952 (
            .O(N__21755),
            .I(N__21735));
    Odrv12 I__3951 (
            .O(N__21752),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    LocalMux I__3950 (
            .O(N__21749),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__3949 (
            .O(N__21744),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv4 I__3948 (
            .O(N__21741),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    LocalMux I__3947 (
            .O(N__21738),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    Odrv12 I__3946 (
            .O(N__21735),
            .I(\this_ppu.M_state_qZ0Z_4 ));
    InMux I__3945 (
            .O(N__21722),
            .I(N__21718));
    InMux I__3944 (
            .O(N__21721),
            .I(N__21715));
    LocalMux I__3943 (
            .O(N__21718),
            .I(N__21711));
    LocalMux I__3942 (
            .O(N__21715),
            .I(N__21706));
    InMux I__3941 (
            .O(N__21714),
            .I(N__21703));
    Span4Mux_v I__3940 (
            .O(N__21711),
            .I(N__21700));
    InMux I__3939 (
            .O(N__21710),
            .I(N__21695));
    InMux I__3938 (
            .O(N__21709),
            .I(N__21695));
    Span4Mux_h I__3937 (
            .O(N__21706),
            .I(N__21690));
    LocalMux I__3936 (
            .O(N__21703),
            .I(N__21690));
    Span4Mux_h I__3935 (
            .O(N__21700),
            .I(N__21685));
    LocalMux I__3934 (
            .O(N__21695),
            .I(N__21685));
    Sp12to4 I__3933 (
            .O(N__21690),
            .I(N__21682));
    Span4Mux_v I__3932 (
            .O(N__21685),
            .I(N__21679));
    Odrv12 I__3931 (
            .O(N__21682),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    Odrv4 I__3930 (
            .O(N__21679),
            .I(\this_ppu.M_state_qZ0Z_10 ));
    CascadeMux I__3929 (
            .O(N__21674),
            .I(\this_ppu.N_835_0_cascade_ ));
    CascadeMux I__3928 (
            .O(N__21671),
            .I(\this_ppu.N_783_cascade_ ));
    InMux I__3927 (
            .O(N__21668),
            .I(N__21665));
    LocalMux I__3926 (
            .O(N__21665),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0 ));
    InMux I__3925 (
            .O(N__21662),
            .I(N__21659));
    LocalMux I__3924 (
            .O(N__21659),
            .I(N__21656));
    Span4Mux_v I__3923 (
            .O(N__21656),
            .I(N__21653));
    Span4Mux_h I__3922 (
            .O(N__21653),
            .I(N__21650));
    Odrv4 I__3921 (
            .O(N__21650),
            .I(\this_ppu.oam_cache.mem_2 ));
    InMux I__3920 (
            .O(N__21647),
            .I(N__21644));
    LocalMux I__3919 (
            .O(N__21644),
            .I(N__21640));
    InMux I__3918 (
            .O(N__21643),
            .I(N__21636));
    Span4Mux_v I__3917 (
            .O(N__21640),
            .I(N__21633));
    InMux I__3916 (
            .O(N__21639),
            .I(N__21630));
    LocalMux I__3915 (
            .O(N__21636),
            .I(\this_ppu.N_60_0 ));
    Odrv4 I__3914 (
            .O(N__21633),
            .I(\this_ppu.N_60_0 ));
    LocalMux I__3913 (
            .O(N__21630),
            .I(\this_ppu.N_60_0 ));
    InMux I__3912 (
            .O(N__21623),
            .I(N__21617));
    CascadeMux I__3911 (
            .O(N__21622),
            .I(N__21614));
    CascadeMux I__3910 (
            .O(N__21621),
            .I(N__21609));
    InMux I__3909 (
            .O(N__21620),
            .I(N__21605));
    LocalMux I__3908 (
            .O(N__21617),
            .I(N__21602));
    InMux I__3907 (
            .O(N__21614),
            .I(N__21595));
    InMux I__3906 (
            .O(N__21613),
            .I(N__21595));
    InMux I__3905 (
            .O(N__21612),
            .I(N__21595));
    InMux I__3904 (
            .O(N__21609),
            .I(N__21591));
    InMux I__3903 (
            .O(N__21608),
            .I(N__21588));
    LocalMux I__3902 (
            .O(N__21605),
            .I(N__21585));
    Span4Mux_v I__3901 (
            .O(N__21602),
            .I(N__21580));
    LocalMux I__3900 (
            .O(N__21595),
            .I(N__21580));
    InMux I__3899 (
            .O(N__21594),
            .I(N__21576));
    LocalMux I__3898 (
            .O(N__21591),
            .I(N__21571));
    LocalMux I__3897 (
            .O(N__21588),
            .I(N__21571));
    Span4Mux_h I__3896 (
            .O(N__21585),
            .I(N__21562));
    Span4Mux_h I__3895 (
            .O(N__21580),
            .I(N__21562));
    InMux I__3894 (
            .O(N__21579),
            .I(N__21559));
    LocalMux I__3893 (
            .O(N__21576),
            .I(N__21554));
    Span4Mux_v I__3892 (
            .O(N__21571),
            .I(N__21554));
    InMux I__3891 (
            .O(N__21570),
            .I(N__21551));
    InMux I__3890 (
            .O(N__21569),
            .I(N__21548));
    InMux I__3889 (
            .O(N__21568),
            .I(N__21543));
    InMux I__3888 (
            .O(N__21567),
            .I(N__21543));
    Sp12to4 I__3887 (
            .O(N__21562),
            .I(N__21538));
    LocalMux I__3886 (
            .O(N__21559),
            .I(N__21538));
    Span4Mux_h I__3885 (
            .O(N__21554),
            .I(N__21535));
    LocalMux I__3884 (
            .O(N__21551),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__3883 (
            .O(N__21548),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    LocalMux I__3882 (
            .O(N__21543),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv12 I__3881 (
            .O(N__21538),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    Odrv4 I__3880 (
            .O(N__21535),
            .I(\this_ppu.M_state_qZ0Z_0 ));
    CascadeMux I__3879 (
            .O(N__21524),
            .I(N__21516));
    InMux I__3878 (
            .O(N__21523),
            .I(N__21507));
    InMux I__3877 (
            .O(N__21522),
            .I(N__21507));
    InMux I__3876 (
            .O(N__21521),
            .I(N__21507));
    InMux I__3875 (
            .O(N__21520),
            .I(N__21507));
    InMux I__3874 (
            .O(N__21519),
            .I(N__21501));
    InMux I__3873 (
            .O(N__21516),
            .I(N__21498));
    LocalMux I__3872 (
            .O(N__21507),
            .I(N__21495));
    InMux I__3871 (
            .O(N__21506),
            .I(N__21492));
    InMux I__3870 (
            .O(N__21505),
            .I(N__21489));
    InMux I__3869 (
            .O(N__21504),
            .I(N__21486));
    LocalMux I__3868 (
            .O(N__21501),
            .I(N__21483));
    LocalMux I__3867 (
            .O(N__21498),
            .I(N__21480));
    Span4Mux_v I__3866 (
            .O(N__21495),
            .I(N__21477));
    LocalMux I__3865 (
            .O(N__21492),
            .I(N__21473));
    LocalMux I__3864 (
            .O(N__21489),
            .I(N__21468));
    LocalMux I__3863 (
            .O(N__21486),
            .I(N__21468));
    Span4Mux_h I__3862 (
            .O(N__21483),
            .I(N__21465));
    Span4Mux_h I__3861 (
            .O(N__21480),
            .I(N__21460));
    Span4Mux_h I__3860 (
            .O(N__21477),
            .I(N__21460));
    InMux I__3859 (
            .O(N__21476),
            .I(N__21457));
    Span4Mux_h I__3858 (
            .O(N__21473),
            .I(N__21454));
    Span4Mux_h I__3857 (
            .O(N__21468),
            .I(N__21449));
    Span4Mux_v I__3856 (
            .O(N__21465),
            .I(N__21449));
    Odrv4 I__3855 (
            .O(N__21460),
            .I(\this_ppu.N_835_0 ));
    LocalMux I__3854 (
            .O(N__21457),
            .I(\this_ppu.N_835_0 ));
    Odrv4 I__3853 (
            .O(N__21454),
            .I(\this_ppu.N_835_0 ));
    Odrv4 I__3852 (
            .O(N__21449),
            .I(\this_ppu.N_835_0 ));
    InMux I__3851 (
            .O(N__21440),
            .I(N__21431));
    InMux I__3850 (
            .O(N__21439),
            .I(N__21428));
    InMux I__3849 (
            .O(N__21438),
            .I(N__21417));
    InMux I__3848 (
            .O(N__21437),
            .I(N__21417));
    InMux I__3847 (
            .O(N__21436),
            .I(N__21417));
    InMux I__3846 (
            .O(N__21435),
            .I(N__21417));
    InMux I__3845 (
            .O(N__21434),
            .I(N__21417));
    LocalMux I__3844 (
            .O(N__21431),
            .I(N__21414));
    LocalMux I__3843 (
            .O(N__21428),
            .I(N__21409));
    LocalMux I__3842 (
            .O(N__21417),
            .I(N__21409));
    Span4Mux_v I__3841 (
            .O(N__21414),
            .I(N__21406));
    Span4Mux_h I__3840 (
            .O(N__21409),
            .I(N__21403));
    Odrv4 I__3839 (
            .O(N__21406),
            .I(\this_ppu.N_807 ));
    Odrv4 I__3838 (
            .O(N__21403),
            .I(\this_ppu.N_807 ));
    CascadeMux I__3837 (
            .O(N__21398),
            .I(N__21395));
    InMux I__3836 (
            .O(N__21395),
            .I(N__21392));
    LocalMux I__3835 (
            .O(N__21392),
            .I(N__21389));
    Span4Mux_h I__3834 (
            .O(N__21389),
            .I(N__21386));
    Odrv4 I__3833 (
            .O(N__21386),
            .I(M_this_scroll_qZ0Z_8));
    CascadeMux I__3832 (
            .O(N__21383),
            .I(N_829_0_cascade_));
    CascadeMux I__3831 (
            .O(N__21380),
            .I(N_58_0_cascade_));
    InMux I__3830 (
            .O(N__21377),
            .I(N__21369));
    InMux I__3829 (
            .O(N__21376),
            .I(N__21366));
    InMux I__3828 (
            .O(N__21375),
            .I(N__21363));
    CascadeMux I__3827 (
            .O(N__21374),
            .I(N__21360));
    InMux I__3826 (
            .O(N__21373),
            .I(N__21356));
    InMux I__3825 (
            .O(N__21372),
            .I(N__21353));
    LocalMux I__3824 (
            .O(N__21369),
            .I(N__21350));
    LocalMux I__3823 (
            .O(N__21366),
            .I(N__21345));
    LocalMux I__3822 (
            .O(N__21363),
            .I(N__21345));
    InMux I__3821 (
            .O(N__21360),
            .I(N__21342));
    CascadeMux I__3820 (
            .O(N__21359),
            .I(N__21338));
    LocalMux I__3819 (
            .O(N__21356),
            .I(N__21335));
    LocalMux I__3818 (
            .O(N__21353),
            .I(N__21332));
    Span4Mux_v I__3817 (
            .O(N__21350),
            .I(N__21327));
    Span4Mux_v I__3816 (
            .O(N__21345),
            .I(N__21327));
    LocalMux I__3815 (
            .O(N__21342),
            .I(N__21324));
    InMux I__3814 (
            .O(N__21341),
            .I(N__21321));
    InMux I__3813 (
            .O(N__21338),
            .I(N__21318));
    Odrv4 I__3812 (
            .O(N__21335),
            .I(\this_ppu.N_97_mux ));
    Odrv4 I__3811 (
            .O(N__21332),
            .I(\this_ppu.N_97_mux ));
    Odrv4 I__3810 (
            .O(N__21327),
            .I(\this_ppu.N_97_mux ));
    Odrv4 I__3809 (
            .O(N__21324),
            .I(\this_ppu.N_97_mux ));
    LocalMux I__3808 (
            .O(N__21321),
            .I(\this_ppu.N_97_mux ));
    LocalMux I__3807 (
            .O(N__21318),
            .I(\this_ppu.N_97_mux ));
    CascadeMux I__3806 (
            .O(N__21305),
            .I(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_ ));
    InMux I__3805 (
            .O(N__21302),
            .I(N__21299));
    LocalMux I__3804 (
            .O(N__21299),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7 ));
    CascadeMux I__3803 (
            .O(N__21296),
            .I(N__21292));
    InMux I__3802 (
            .O(N__21295),
            .I(N__21289));
    InMux I__3801 (
            .O(N__21292),
            .I(N__21286));
    LocalMux I__3800 (
            .O(N__21289),
            .I(N__21283));
    LocalMux I__3799 (
            .O(N__21286),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_2 ));
    Odrv4 I__3798 (
            .O(N__21283),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_2 ));
    CascadeMux I__3797 (
            .O(N__21278),
            .I(N__21275));
    InMux I__3796 (
            .O(N__21275),
            .I(N__21271));
    InMux I__3795 (
            .O(N__21274),
            .I(N__21268));
    LocalMux I__3794 (
            .O(N__21271),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_1 ));
    LocalMux I__3793 (
            .O(N__21268),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_1 ));
    CascadeMux I__3792 (
            .O(N__21263),
            .I(N__21259));
    CascadeMux I__3791 (
            .O(N__21262),
            .I(N__21256));
    InMux I__3790 (
            .O(N__21259),
            .I(N__21253));
    InMux I__3789 (
            .O(N__21256),
            .I(N__21250));
    LocalMux I__3788 (
            .O(N__21253),
            .I(N__21247));
    LocalMux I__3787 (
            .O(N__21250),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_7 ));
    Odrv4 I__3786 (
            .O(N__21247),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_7 ));
    InMux I__3785 (
            .O(N__21242),
            .I(N__21239));
    LocalMux I__3784 (
            .O(N__21239),
            .I(\this_ppu.m9_0_a2_4 ));
    InMux I__3783 (
            .O(N__21236),
            .I(N__21232));
    CascadeMux I__3782 (
            .O(N__21235),
            .I(N__21228));
    LocalMux I__3781 (
            .O(N__21232),
            .I(N__21225));
    InMux I__3780 (
            .O(N__21231),
            .I(N__21222));
    InMux I__3779 (
            .O(N__21228),
            .I(N__21219));
    Span4Mux_v I__3778 (
            .O(N__21225),
            .I(N__21214));
    LocalMux I__3777 (
            .O(N__21222),
            .I(N__21214));
    LocalMux I__3776 (
            .O(N__21219),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_0 ));
    Odrv4 I__3775 (
            .O(N__21214),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_0 ));
    InMux I__3774 (
            .O(N__21209),
            .I(N__21206));
    LocalMux I__3773 (
            .O(N__21206),
            .I(N__21203));
    Span4Mux_v I__3772 (
            .O(N__21203),
            .I(N__21200));
    Odrv4 I__3771 (
            .O(N__21200),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_axb_0 ));
    InMux I__3770 (
            .O(N__21197),
            .I(N__21194));
    LocalMux I__3769 (
            .O(N__21194),
            .I(\this_ppu.un1_M_surface_x_q_c2 ));
    InMux I__3768 (
            .O(N__21191),
            .I(N__21183));
    InMux I__3767 (
            .O(N__21190),
            .I(N__21183));
    InMux I__3766 (
            .O(N__21189),
            .I(N__21180));
    InMux I__3765 (
            .O(N__21188),
            .I(N__21177));
    LocalMux I__3764 (
            .O(N__21183),
            .I(\this_ppu.M_oam_curr_dZ0Z25 ));
    LocalMux I__3763 (
            .O(N__21180),
            .I(\this_ppu.M_oam_curr_dZ0Z25 ));
    LocalMux I__3762 (
            .O(N__21177),
            .I(\this_ppu.M_oam_curr_dZ0Z25 ));
    InMux I__3761 (
            .O(N__21170),
            .I(N__21167));
    LocalMux I__3760 (
            .O(N__21167),
            .I(N__21160));
    CascadeMux I__3759 (
            .O(N__21166),
            .I(N__21157));
    InMux I__3758 (
            .O(N__21165),
            .I(N__21152));
    InMux I__3757 (
            .O(N__21164),
            .I(N__21149));
    InMux I__3756 (
            .O(N__21163),
            .I(N__21146));
    Span4Mux_v I__3755 (
            .O(N__21160),
            .I(N__21143));
    InMux I__3754 (
            .O(N__21157),
            .I(N__21140));
    InMux I__3753 (
            .O(N__21156),
            .I(N__21135));
    InMux I__3752 (
            .O(N__21155),
            .I(N__21135));
    LocalMux I__3751 (
            .O(N__21152),
            .I(N__21130));
    LocalMux I__3750 (
            .O(N__21149),
            .I(N__21130));
    LocalMux I__3749 (
            .O(N__21146),
            .I(N__21127));
    Odrv4 I__3748 (
            .O(N__21143),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__3747 (
            .O(N__21140),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    LocalMux I__3746 (
            .O(N__21135),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__3745 (
            .O(N__21130),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    Odrv4 I__3744 (
            .O(N__21127),
            .I(\this_ppu.M_state_qZ0Z_7 ));
    CascadeMux I__3743 (
            .O(N__21116),
            .I(N__21109));
    CascadeMux I__3742 (
            .O(N__21115),
            .I(N__21106));
    InMux I__3741 (
            .O(N__21114),
            .I(N__21103));
    InMux I__3740 (
            .O(N__21113),
            .I(N__21100));
    InMux I__3739 (
            .O(N__21112),
            .I(N__21092));
    InMux I__3738 (
            .O(N__21109),
            .I(N__21092));
    InMux I__3737 (
            .O(N__21106),
            .I(N__21092));
    LocalMux I__3736 (
            .O(N__21103),
            .I(N__21086));
    LocalMux I__3735 (
            .O(N__21100),
            .I(N__21086));
    InMux I__3734 (
            .O(N__21099),
            .I(N__21083));
    LocalMux I__3733 (
            .O(N__21092),
            .I(N__21080));
    InMux I__3732 (
            .O(N__21091),
            .I(N__21077));
    Span4Mux_v I__3731 (
            .O(N__21086),
            .I(N__21074));
    LocalMux I__3730 (
            .O(N__21083),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv4 I__3729 (
            .O(N__21080),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    LocalMux I__3728 (
            .O(N__21077),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    Odrv4 I__3727 (
            .O(N__21074),
            .I(\this_ppu.M_state_qZ0Z_9 ));
    CascadeMux I__3726 (
            .O(N__21065),
            .I(\this_ppu.un1_M_surface_x_q_c1_cascade_ ));
    CascadeMux I__3725 (
            .O(N__21062),
            .I(N__21059));
    InMux I__3724 (
            .O(N__21059),
            .I(N__21056));
    LocalMux I__3723 (
            .O(N__21056),
            .I(N__21053));
    Odrv4 I__3722 (
            .O(N__21053),
            .I(M_this_scroll_qZ0Z_10));
    InMux I__3721 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__3720 (
            .O(N__21047),
            .I(N__21044));
    Odrv4 I__3719 (
            .O(N__21044),
            .I(M_this_scroll_qZ0Z_11));
    InMux I__3718 (
            .O(N__21041),
            .I(N__21038));
    LocalMux I__3717 (
            .O(N__21038),
            .I(M_this_scroll_qZ0Z_13));
    InMux I__3716 (
            .O(N__21035),
            .I(N__21032));
    LocalMux I__3715 (
            .O(N__21032),
            .I(N__21029));
    Span4Mux_v I__3714 (
            .O(N__21029),
            .I(N__21026));
    Odrv4 I__3713 (
            .O(N__21026),
            .I(M_this_scroll_qZ0Z_14));
    CascadeMux I__3712 (
            .O(N__21023),
            .I(\this_ppu.N_798_0_cascade_ ));
    CascadeMux I__3711 (
            .O(N__21020),
            .I(N__21017));
    InMux I__3710 (
            .O(N__21017),
            .I(N__21014));
    LocalMux I__3709 (
            .O(N__21014),
            .I(\this_ppu.un1_M_surface_x_q_c3 ));
    CascadeMux I__3708 (
            .O(N__21011),
            .I(\this_ppu.un1_M_surface_x_q_c3_cascade_ ));
    InMux I__3707 (
            .O(N__21008),
            .I(N__21005));
    LocalMux I__3706 (
            .O(N__21005),
            .I(\this_ppu.N_798_0 ));
    CascadeMux I__3705 (
            .O(N__21002),
            .I(\this_ppu.un1_M_surface_x_q_c2_cascade_ ));
    CascadeMux I__3704 (
            .O(N__20999),
            .I(\this_ppu.un1_M_surface_x_q_c5_cascade_ ));
    InMux I__3703 (
            .O(N__20996),
            .I(N__20993));
    LocalMux I__3702 (
            .O(N__20993),
            .I(N__20989));
    InMux I__3701 (
            .O(N__20992),
            .I(N__20986));
    Odrv4 I__3700 (
            .O(N__20989),
            .I(\this_ppu.N_800 ));
    LocalMux I__3699 (
            .O(N__20986),
            .I(\this_ppu.N_800 ));
    CascadeMux I__3698 (
            .O(N__20981),
            .I(\this_ppu.N_800_cascade_ ));
    InMux I__3697 (
            .O(N__20978),
            .I(N__20972));
    CascadeMux I__3696 (
            .O(N__20977),
            .I(N__20968));
    InMux I__3695 (
            .O(N__20976),
            .I(N__20965));
    InMux I__3694 (
            .O(N__20975),
            .I(N__20962));
    LocalMux I__3693 (
            .O(N__20972),
            .I(N__20959));
    InMux I__3692 (
            .O(N__20971),
            .I(N__20956));
    InMux I__3691 (
            .O(N__20968),
            .I(N__20953));
    LocalMux I__3690 (
            .O(N__20965),
            .I(N__20948));
    LocalMux I__3689 (
            .O(N__20962),
            .I(N__20948));
    Span4Mux_v I__3688 (
            .O(N__20959),
            .I(N__20941));
    LocalMux I__3687 (
            .O(N__20956),
            .I(N__20941));
    LocalMux I__3686 (
            .O(N__20953),
            .I(N__20941));
    Span4Mux_h I__3685 (
            .O(N__20948),
            .I(N__20938));
    Span4Mux_v I__3684 (
            .O(N__20941),
            .I(N__20935));
    Odrv4 I__3683 (
            .O(N__20938),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    Odrv4 I__3682 (
            .O(N__20935),
            .I(\this_ppu.M_state_qZ0Z_11 ));
    CEMux I__3681 (
            .O(N__20930),
            .I(N__20927));
    LocalMux I__3680 (
            .O(N__20927),
            .I(N__20924));
    Span4Mux_v I__3679 (
            .O(N__20924),
            .I(N__20921));
    Span4Mux_h I__3678 (
            .O(N__20921),
            .I(N__20918));
    Odrv4 I__3677 (
            .O(N__20918),
            .I(N_18));
    CascadeMux I__3676 (
            .O(N__20915),
            .I(\this_ppu.un3_M_screen_y_d_0_c4_cascade_ ));
    CascadeMux I__3675 (
            .O(N__20912),
            .I(N__20909));
    InMux I__3674 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__3673 (
            .O(N__20906),
            .I(N__20903));
    Span4Mux_h I__3672 (
            .O(N__20903),
            .I(N__20900));
    Odrv4 I__3671 (
            .O(N__20900),
            .I(\this_ppu.N_802 ));
    InMux I__3670 (
            .O(N__20897),
            .I(N__20894));
    LocalMux I__3669 (
            .O(N__20894),
            .I(N__20891));
    Span12Mux_h I__3668 (
            .O(N__20891),
            .I(N__20888));
    Span12Mux_v I__3667 (
            .O(N__20888),
            .I(N__20885));
    Odrv12 I__3666 (
            .O(N__20885),
            .I(\this_spr_ram.mem_out_bus7_3 ));
    InMux I__3665 (
            .O(N__20882),
            .I(N__20879));
    LocalMux I__3664 (
            .O(N__20879),
            .I(N__20876));
    Span12Mux_v I__3663 (
            .O(N__20876),
            .I(N__20873));
    Span12Mux_h I__3662 (
            .O(N__20873),
            .I(N__20870));
    Odrv12 I__3661 (
            .O(N__20870),
            .I(\this_spr_ram.mem_out_bus3_3 ));
    InMux I__3660 (
            .O(N__20867),
            .I(N__20860));
    InMux I__3659 (
            .O(N__20866),
            .I(N__20853));
    InMux I__3658 (
            .O(N__20865),
            .I(N__20853));
    InMux I__3657 (
            .O(N__20864),
            .I(N__20853));
    InMux I__3656 (
            .O(N__20863),
            .I(N__20849));
    LocalMux I__3655 (
            .O(N__20860),
            .I(N__20844));
    LocalMux I__3654 (
            .O(N__20853),
            .I(N__20844));
    InMux I__3653 (
            .O(N__20852),
            .I(N__20841));
    LocalMux I__3652 (
            .O(N__20849),
            .I(N__20831));
    Span4Mux_v I__3651 (
            .O(N__20844),
            .I(N__20831));
    LocalMux I__3650 (
            .O(N__20841),
            .I(N__20831));
    InMux I__3649 (
            .O(N__20840),
            .I(N__20819));
    InMux I__3648 (
            .O(N__20839),
            .I(N__20819));
    InMux I__3647 (
            .O(N__20838),
            .I(N__20816));
    Span4Mux_v I__3646 (
            .O(N__20831),
            .I(N__20813));
    InMux I__3645 (
            .O(N__20830),
            .I(N__20806));
    InMux I__3644 (
            .O(N__20829),
            .I(N__20806));
    InMux I__3643 (
            .O(N__20828),
            .I(N__20806));
    InMux I__3642 (
            .O(N__20827),
            .I(N__20801));
    InMux I__3641 (
            .O(N__20826),
            .I(N__20801));
    InMux I__3640 (
            .O(N__20825),
            .I(N__20798));
    InMux I__3639 (
            .O(N__20824),
            .I(N__20795));
    LocalMux I__3638 (
            .O(N__20819),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__3637 (
            .O(N__20816),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    Odrv4 I__3636 (
            .O(N__20813),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__3635 (
            .O(N__20806),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__3634 (
            .O(N__20801),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__3633 (
            .O(N__20798),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    LocalMux I__3632 (
            .O(N__20795),
            .I(\this_spr_ram.mem_radregZ0Z_13 ));
    InMux I__3631 (
            .O(N__20780),
            .I(N__20777));
    LocalMux I__3630 (
            .O(N__20777),
            .I(N__20774));
    Odrv4 I__3629 (
            .O(N__20774),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ));
    InMux I__3628 (
            .O(N__20771),
            .I(N__20764));
    InMux I__3627 (
            .O(N__20770),
            .I(N__20761));
    InMux I__3626 (
            .O(N__20769),
            .I(N__20756));
    InMux I__3625 (
            .O(N__20768),
            .I(N__20756));
    InMux I__3624 (
            .O(N__20767),
            .I(N__20753));
    LocalMux I__3623 (
            .O(N__20764),
            .I(N__20750));
    LocalMux I__3622 (
            .O(N__20761),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__3621 (
            .O(N__20756),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    LocalMux I__3620 (
            .O(N__20753),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    Odrv12 I__3619 (
            .O(N__20750),
            .I(\this_ppu.M_state_qZ0Z_5 ));
    CascadeMux I__3618 (
            .O(N__20741),
            .I(N__20738));
    InMux I__3617 (
            .O(N__20738),
            .I(N__20734));
    InMux I__3616 (
            .O(N__20737),
            .I(N__20731));
    LocalMux I__3615 (
            .O(N__20734),
            .I(N__20726));
    LocalMux I__3614 (
            .O(N__20731),
            .I(N__20726));
    Span4Mux_v I__3613 (
            .O(N__20726),
            .I(N__20723));
    Span4Mux_h I__3612 (
            .O(N__20723),
            .I(N__20720));
    Span4Mux_v I__3611 (
            .O(N__20720),
            .I(N__20717));
    Odrv4 I__3610 (
            .O(N__20717),
            .I(\this_ppu.N_796_0 ));
    InMux I__3609 (
            .O(N__20714),
            .I(N__20711));
    LocalMux I__3608 (
            .O(N__20711),
            .I(\this_ppu.M_state_qZ0Z_8 ));
    CascadeMux I__3607 (
            .O(N__20708),
            .I(\this_ppu.un1_M_surface_x_q_c6_cascade_ ));
    InMux I__3606 (
            .O(N__20705),
            .I(N__20702));
    LocalMux I__3605 (
            .O(N__20702),
            .I(N__20699));
    Span12Mux_v I__3604 (
            .O(N__20699),
            .I(N__20696));
    Span12Mux_h I__3603 (
            .O(N__20696),
            .I(N__20693));
    Odrv12 I__3602 (
            .O(N__20693),
            .I(M_this_map_ram_read_data_7));
    InMux I__3601 (
            .O(N__20690),
            .I(N__20687));
    LocalMux I__3600 (
            .O(N__20687),
            .I(N__20684));
    Odrv12 I__3599 (
            .O(N__20684),
            .I(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ));
    InMux I__3598 (
            .O(N__20681),
            .I(N__20678));
    LocalMux I__3597 (
            .O(N__20678),
            .I(N__20675));
    Span4Mux_h I__3596 (
            .O(N__20675),
            .I(N__20672));
    Odrv4 I__3595 (
            .O(N__20672),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_3 ));
    InMux I__3594 (
            .O(N__20669),
            .I(N__20666));
    LocalMux I__3593 (
            .O(N__20666),
            .I(N__20663));
    Span4Mux_h I__3592 (
            .O(N__20663),
            .I(N__20660));
    Span4Mux_h I__3591 (
            .O(N__20660),
            .I(N__20657));
    Sp12to4 I__3590 (
            .O(N__20657),
            .I(N__20654));
    Span12Mux_v I__3589 (
            .O(N__20654),
            .I(N__20651));
    Odrv12 I__3588 (
            .O(N__20651),
            .I(M_this_map_ram_read_data_3));
    CascadeMux I__3587 (
            .O(N__20648),
            .I(N__20644));
    CascadeMux I__3586 (
            .O(N__20647),
            .I(N__20641));
    InMux I__3585 (
            .O(N__20644),
            .I(N__20634));
    InMux I__3584 (
            .O(N__20641),
            .I(N__20631));
    CascadeMux I__3583 (
            .O(N__20640),
            .I(N__20628));
    CascadeMux I__3582 (
            .O(N__20639),
            .I(N__20624));
    CascadeMux I__3581 (
            .O(N__20638),
            .I(N__20616));
    CascadeMux I__3580 (
            .O(N__20637),
            .I(N__20613));
    LocalMux I__3579 (
            .O(N__20634),
            .I(N__20607));
    LocalMux I__3578 (
            .O(N__20631),
            .I(N__20607));
    InMux I__3577 (
            .O(N__20628),
            .I(N__20604));
    CascadeMux I__3576 (
            .O(N__20627),
            .I(N__20601));
    InMux I__3575 (
            .O(N__20624),
            .I(N__20598));
    CascadeMux I__3574 (
            .O(N__20623),
            .I(N__20595));
    CascadeMux I__3573 (
            .O(N__20622),
            .I(N__20592));
    CascadeMux I__3572 (
            .O(N__20621),
            .I(N__20589));
    CascadeMux I__3571 (
            .O(N__20620),
            .I(N__20585));
    CascadeMux I__3570 (
            .O(N__20619),
            .I(N__20582));
    InMux I__3569 (
            .O(N__20616),
            .I(N__20577));
    InMux I__3568 (
            .O(N__20613),
            .I(N__20574));
    CascadeMux I__3567 (
            .O(N__20612),
            .I(N__20571));
    Span4Mux_s2_v I__3566 (
            .O(N__20607),
            .I(N__20566));
    LocalMux I__3565 (
            .O(N__20604),
            .I(N__20566));
    InMux I__3564 (
            .O(N__20601),
            .I(N__20563));
    LocalMux I__3563 (
            .O(N__20598),
            .I(N__20560));
    InMux I__3562 (
            .O(N__20595),
            .I(N__20557));
    InMux I__3561 (
            .O(N__20592),
            .I(N__20554));
    InMux I__3560 (
            .O(N__20589),
            .I(N__20551));
    CascadeMux I__3559 (
            .O(N__20588),
            .I(N__20548));
    InMux I__3558 (
            .O(N__20585),
            .I(N__20545));
    InMux I__3557 (
            .O(N__20582),
            .I(N__20542));
    CascadeMux I__3556 (
            .O(N__20581),
            .I(N__20539));
    CascadeMux I__3555 (
            .O(N__20580),
            .I(N__20536));
    LocalMux I__3554 (
            .O(N__20577),
            .I(N__20533));
    LocalMux I__3553 (
            .O(N__20574),
            .I(N__20530));
    InMux I__3552 (
            .O(N__20571),
            .I(N__20527));
    Span4Mux_v I__3551 (
            .O(N__20566),
            .I(N__20522));
    LocalMux I__3550 (
            .O(N__20563),
            .I(N__20522));
    Span4Mux_v I__3549 (
            .O(N__20560),
            .I(N__20517));
    LocalMux I__3548 (
            .O(N__20557),
            .I(N__20517));
    LocalMux I__3547 (
            .O(N__20554),
            .I(N__20514));
    LocalMux I__3546 (
            .O(N__20551),
            .I(N__20511));
    InMux I__3545 (
            .O(N__20548),
            .I(N__20508));
    LocalMux I__3544 (
            .O(N__20545),
            .I(N__20503));
    LocalMux I__3543 (
            .O(N__20542),
            .I(N__20503));
    InMux I__3542 (
            .O(N__20539),
            .I(N__20500));
    InMux I__3541 (
            .O(N__20536),
            .I(N__20497));
    Span4Mux_v I__3540 (
            .O(N__20533),
            .I(N__20492));
    Span4Mux_v I__3539 (
            .O(N__20530),
            .I(N__20492));
    LocalMux I__3538 (
            .O(N__20527),
            .I(N__20489));
    Span4Mux_h I__3537 (
            .O(N__20522),
            .I(N__20486));
    Span4Mux_v I__3536 (
            .O(N__20517),
            .I(N__20477));
    Span4Mux_v I__3535 (
            .O(N__20514),
            .I(N__20477));
    Span4Mux_v I__3534 (
            .O(N__20511),
            .I(N__20477));
    LocalMux I__3533 (
            .O(N__20508),
            .I(N__20477));
    Span4Mux_s2_v I__3532 (
            .O(N__20503),
            .I(N__20472));
    LocalMux I__3531 (
            .O(N__20500),
            .I(N__20472));
    LocalMux I__3530 (
            .O(N__20497),
            .I(N__20469));
    Sp12to4 I__3529 (
            .O(N__20492),
            .I(N__20464));
    Span12Mux_s8_h I__3528 (
            .O(N__20489),
            .I(N__20464));
    Span4Mux_v I__3527 (
            .O(N__20486),
            .I(N__20459));
    Span4Mux_h I__3526 (
            .O(N__20477),
            .I(N__20459));
    Span4Mux_v I__3525 (
            .O(N__20472),
            .I(N__20454));
    Span4Mux_h I__3524 (
            .O(N__20469),
            .I(N__20454));
    Span12Mux_v I__3523 (
            .O(N__20464),
            .I(N__20449));
    Sp12to4 I__3522 (
            .O(N__20459),
            .I(N__20449));
    Span4Mux_h I__3521 (
            .O(N__20454),
            .I(N__20446));
    Odrv12 I__3520 (
            .O(N__20449),
            .I(M_this_ppu_spr_addr_9));
    Odrv4 I__3519 (
            .O(N__20446),
            .I(M_this_ppu_spr_addr_9));
    InMux I__3518 (
            .O(N__20441),
            .I(N__20438));
    LocalMux I__3517 (
            .O(N__20438),
            .I(N__20435));
    Span4Mux_h I__3516 (
            .O(N__20435),
            .I(N__20432));
    Odrv4 I__3515 (
            .O(N__20432),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_4 ));
    InMux I__3514 (
            .O(N__20429),
            .I(N__20426));
    LocalMux I__3513 (
            .O(N__20426),
            .I(N__20423));
    Span4Mux_v I__3512 (
            .O(N__20423),
            .I(N__20420));
    Span4Mux_v I__3511 (
            .O(N__20420),
            .I(N__20417));
    Sp12to4 I__3510 (
            .O(N__20417),
            .I(N__20414));
    Span12Mux_h I__3509 (
            .O(N__20414),
            .I(N__20411));
    Span12Mux_v I__3508 (
            .O(N__20411),
            .I(N__20408));
    Odrv12 I__3507 (
            .O(N__20408),
            .I(M_this_map_ram_read_data_4));
    CascadeMux I__3506 (
            .O(N__20405),
            .I(N__20402));
    InMux I__3505 (
            .O(N__20402),
            .I(N__20397));
    CascadeMux I__3504 (
            .O(N__20401),
            .I(N__20394));
    CascadeMux I__3503 (
            .O(N__20400),
            .I(N__20390));
    LocalMux I__3502 (
            .O(N__20397),
            .I(N__20386));
    InMux I__3501 (
            .O(N__20394),
            .I(N__20383));
    CascadeMux I__3500 (
            .O(N__20393),
            .I(N__20380));
    InMux I__3499 (
            .O(N__20390),
            .I(N__20374));
    CascadeMux I__3498 (
            .O(N__20389),
            .I(N__20371));
    Span4Mux_s2_v I__3497 (
            .O(N__20386),
            .I(N__20366));
    LocalMux I__3496 (
            .O(N__20383),
            .I(N__20366));
    InMux I__3495 (
            .O(N__20380),
            .I(N__20363));
    CascadeMux I__3494 (
            .O(N__20379),
            .I(N__20360));
    CascadeMux I__3493 (
            .O(N__20378),
            .I(N__20356));
    CascadeMux I__3492 (
            .O(N__20377),
            .I(N__20353));
    LocalMux I__3491 (
            .O(N__20374),
            .I(N__20347));
    InMux I__3490 (
            .O(N__20371),
            .I(N__20344));
    Span4Mux_h I__3489 (
            .O(N__20366),
            .I(N__20338));
    LocalMux I__3488 (
            .O(N__20363),
            .I(N__20338));
    InMux I__3487 (
            .O(N__20360),
            .I(N__20335));
    CascadeMux I__3486 (
            .O(N__20359),
            .I(N__20332));
    InMux I__3485 (
            .O(N__20356),
            .I(N__20329));
    InMux I__3484 (
            .O(N__20353),
            .I(N__20326));
    CascadeMux I__3483 (
            .O(N__20352),
            .I(N__20323));
    CascadeMux I__3482 (
            .O(N__20351),
            .I(N__20319));
    CascadeMux I__3481 (
            .O(N__20350),
            .I(N__20316));
    Span4Mux_h I__3480 (
            .O(N__20347),
            .I(N__20309));
    LocalMux I__3479 (
            .O(N__20344),
            .I(N__20309));
    CascadeMux I__3478 (
            .O(N__20343),
            .I(N__20306));
    Span4Mux_v I__3477 (
            .O(N__20338),
            .I(N__20301));
    LocalMux I__3476 (
            .O(N__20335),
            .I(N__20301));
    InMux I__3475 (
            .O(N__20332),
            .I(N__20298));
    LocalMux I__3474 (
            .O(N__20329),
            .I(N__20295));
    LocalMux I__3473 (
            .O(N__20326),
            .I(N__20292));
    InMux I__3472 (
            .O(N__20323),
            .I(N__20289));
    CascadeMux I__3471 (
            .O(N__20322),
            .I(N__20286));
    InMux I__3470 (
            .O(N__20319),
            .I(N__20283));
    InMux I__3469 (
            .O(N__20316),
            .I(N__20280));
    CascadeMux I__3468 (
            .O(N__20315),
            .I(N__20277));
    CascadeMux I__3467 (
            .O(N__20314),
            .I(N__20274));
    Span4Mux_v I__3466 (
            .O(N__20309),
            .I(N__20271));
    InMux I__3465 (
            .O(N__20306),
            .I(N__20268));
    Span4Mux_h I__3464 (
            .O(N__20301),
            .I(N__20263));
    LocalMux I__3463 (
            .O(N__20298),
            .I(N__20263));
    Span4Mux_v I__3462 (
            .O(N__20295),
            .I(N__20256));
    Span4Mux_h I__3461 (
            .O(N__20292),
            .I(N__20256));
    LocalMux I__3460 (
            .O(N__20289),
            .I(N__20256));
    InMux I__3459 (
            .O(N__20286),
            .I(N__20253));
    LocalMux I__3458 (
            .O(N__20283),
            .I(N__20248));
    LocalMux I__3457 (
            .O(N__20280),
            .I(N__20248));
    InMux I__3456 (
            .O(N__20277),
            .I(N__20245));
    InMux I__3455 (
            .O(N__20274),
            .I(N__20242));
    Sp12to4 I__3454 (
            .O(N__20271),
            .I(N__20237));
    LocalMux I__3453 (
            .O(N__20268),
            .I(N__20237));
    Span4Mux_v I__3452 (
            .O(N__20263),
            .I(N__20230));
    Span4Mux_v I__3451 (
            .O(N__20256),
            .I(N__20230));
    LocalMux I__3450 (
            .O(N__20253),
            .I(N__20230));
    Span4Mux_s2_v I__3449 (
            .O(N__20248),
            .I(N__20225));
    LocalMux I__3448 (
            .O(N__20245),
            .I(N__20225));
    LocalMux I__3447 (
            .O(N__20242),
            .I(N__20222));
    Span12Mux_h I__3446 (
            .O(N__20237),
            .I(N__20219));
    Sp12to4 I__3445 (
            .O(N__20230),
            .I(N__20216));
    Span4Mux_v I__3444 (
            .O(N__20225),
            .I(N__20211));
    Span4Mux_h I__3443 (
            .O(N__20222),
            .I(N__20211));
    Span12Mux_v I__3442 (
            .O(N__20219),
            .I(N__20206));
    Span12Mux_h I__3441 (
            .O(N__20216),
            .I(N__20206));
    Span4Mux_h I__3440 (
            .O(N__20211),
            .I(N__20203));
    Odrv12 I__3439 (
            .O(N__20206),
            .I(M_this_ppu_spr_addr_10));
    Odrv4 I__3438 (
            .O(N__20203),
            .I(M_this_ppu_spr_addr_10));
    CascadeMux I__3437 (
            .O(N__20198),
            .I(N__20193));
    CascadeMux I__3436 (
            .O(N__20197),
            .I(N__20189));
    CascadeMux I__3435 (
            .O(N__20196),
            .I(N__20186));
    InMux I__3434 (
            .O(N__20193),
            .I(N__20182));
    CascadeMux I__3433 (
            .O(N__20192),
            .I(N__20179));
    InMux I__3432 (
            .O(N__20189),
            .I(N__20173));
    InMux I__3431 (
            .O(N__20186),
            .I(N__20170));
    CascadeMux I__3430 (
            .O(N__20185),
            .I(N__20166));
    LocalMux I__3429 (
            .O(N__20182),
            .I(N__20162));
    InMux I__3428 (
            .O(N__20179),
            .I(N__20159));
    CascadeMux I__3427 (
            .O(N__20178),
            .I(N__20156));
    CascadeMux I__3426 (
            .O(N__20177),
            .I(N__20152));
    CascadeMux I__3425 (
            .O(N__20176),
            .I(N__20149));
    LocalMux I__3424 (
            .O(N__20173),
            .I(N__20140));
    LocalMux I__3423 (
            .O(N__20170),
            .I(N__20140));
    CascadeMux I__3422 (
            .O(N__20169),
            .I(N__20137));
    InMux I__3421 (
            .O(N__20166),
            .I(N__20134));
    CascadeMux I__3420 (
            .O(N__20165),
            .I(N__20131));
    Span4Mux_v I__3419 (
            .O(N__20162),
            .I(N__20126));
    LocalMux I__3418 (
            .O(N__20159),
            .I(N__20126));
    InMux I__3417 (
            .O(N__20156),
            .I(N__20123));
    CascadeMux I__3416 (
            .O(N__20155),
            .I(N__20120));
    InMux I__3415 (
            .O(N__20152),
            .I(N__20116));
    InMux I__3414 (
            .O(N__20149),
            .I(N__20113));
    CascadeMux I__3413 (
            .O(N__20148),
            .I(N__20110));
    CascadeMux I__3412 (
            .O(N__20147),
            .I(N__20107));
    CascadeMux I__3411 (
            .O(N__20146),
            .I(N__20104));
    CascadeMux I__3410 (
            .O(N__20145),
            .I(N__20101));
    Span4Mux_v I__3409 (
            .O(N__20140),
            .I(N__20098));
    InMux I__3408 (
            .O(N__20137),
            .I(N__20095));
    LocalMux I__3407 (
            .O(N__20134),
            .I(N__20092));
    InMux I__3406 (
            .O(N__20131),
            .I(N__20089));
    Span4Mux_h I__3405 (
            .O(N__20126),
            .I(N__20084));
    LocalMux I__3404 (
            .O(N__20123),
            .I(N__20084));
    InMux I__3403 (
            .O(N__20120),
            .I(N__20081));
    CascadeMux I__3402 (
            .O(N__20119),
            .I(N__20078));
    LocalMux I__3401 (
            .O(N__20116),
            .I(N__20073));
    LocalMux I__3400 (
            .O(N__20113),
            .I(N__20073));
    InMux I__3399 (
            .O(N__20110),
            .I(N__20070));
    InMux I__3398 (
            .O(N__20107),
            .I(N__20067));
    InMux I__3397 (
            .O(N__20104),
            .I(N__20064));
    InMux I__3396 (
            .O(N__20101),
            .I(N__20061));
    Span4Mux_h I__3395 (
            .O(N__20098),
            .I(N__20058));
    LocalMux I__3394 (
            .O(N__20095),
            .I(N__20055));
    Span4Mux_v I__3393 (
            .O(N__20092),
            .I(N__20046));
    LocalMux I__3392 (
            .O(N__20089),
            .I(N__20046));
    Span4Mux_v I__3391 (
            .O(N__20084),
            .I(N__20046));
    LocalMux I__3390 (
            .O(N__20081),
            .I(N__20046));
    InMux I__3389 (
            .O(N__20078),
            .I(N__20043));
    Span4Mux_s2_v I__3388 (
            .O(N__20073),
            .I(N__20038));
    LocalMux I__3387 (
            .O(N__20070),
            .I(N__20038));
    LocalMux I__3386 (
            .O(N__20067),
            .I(N__20035));
    LocalMux I__3385 (
            .O(N__20064),
            .I(N__20030));
    LocalMux I__3384 (
            .O(N__20061),
            .I(N__20030));
    Sp12to4 I__3383 (
            .O(N__20058),
            .I(N__20025));
    Span12Mux_h I__3382 (
            .O(N__20055),
            .I(N__20025));
    Span4Mux_v I__3381 (
            .O(N__20046),
            .I(N__20022));
    LocalMux I__3380 (
            .O(N__20043),
            .I(N__20019));
    Span4Mux_v I__3379 (
            .O(N__20038),
            .I(N__20014));
    Span4Mux_h I__3378 (
            .O(N__20035),
            .I(N__20014));
    Span12Mux_s10_v I__3377 (
            .O(N__20030),
            .I(N__20005));
    Span12Mux_v I__3376 (
            .O(N__20025),
            .I(N__20005));
    Sp12to4 I__3375 (
            .O(N__20022),
            .I(N__20005));
    Span12Mux_s7_h I__3374 (
            .O(N__20019),
            .I(N__20005));
    Span4Mux_h I__3373 (
            .O(N__20014),
            .I(N__20002));
    Odrv12 I__3372 (
            .O(N__20005),
            .I(M_this_ppu_spr_addr_0));
    Odrv4 I__3371 (
            .O(N__20002),
            .I(M_this_ppu_spr_addr_0));
    InMux I__3370 (
            .O(N__19997),
            .I(N__19994));
    LocalMux I__3369 (
            .O(N__19994),
            .I(N__19991));
    Span12Mux_h I__3368 (
            .O(N__19991),
            .I(N__19988));
    Span12Mux_v I__3367 (
            .O(N__19988),
            .I(N__19985));
    Odrv12 I__3366 (
            .O(N__19985),
            .I(\this_spr_ram.mem_out_bus6_3 ));
    InMux I__3365 (
            .O(N__19982),
            .I(N__19979));
    LocalMux I__3364 (
            .O(N__19979),
            .I(N__19976));
    Span12Mux_v I__3363 (
            .O(N__19976),
            .I(N__19973));
    Span12Mux_h I__3362 (
            .O(N__19973),
            .I(N__19970));
    Odrv12 I__3361 (
            .O(N__19970),
            .I(\this_spr_ram.mem_out_bus2_3 ));
    InMux I__3360 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__3359 (
            .O(N__19964),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ));
    InMux I__3358 (
            .O(N__19961),
            .I(N__19958));
    LocalMux I__3357 (
            .O(N__19958),
            .I(N__19955));
    Span4Mux_h I__3356 (
            .O(N__19955),
            .I(N__19952));
    Odrv4 I__3355 (
            .O(N__19952),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_5 ));
    InMux I__3354 (
            .O(N__19949),
            .I(N__19946));
    LocalMux I__3353 (
            .O(N__19946),
            .I(N__19943));
    Span4Mux_h I__3352 (
            .O(N__19943),
            .I(N__19940));
    Sp12to4 I__3351 (
            .O(N__19940),
            .I(N__19937));
    Span12Mux_v I__3350 (
            .O(N__19937),
            .I(N__19934));
    Span12Mux_h I__3349 (
            .O(N__19934),
            .I(N__19931));
    Odrv12 I__3348 (
            .O(N__19931),
            .I(M_this_map_ram_read_data_5));
    CascadeMux I__3347 (
            .O(N__19928),
            .I(N__19922));
    InMux I__3346 (
            .O(N__19927),
            .I(N__19919));
    InMux I__3345 (
            .O(N__19926),
            .I(N__19916));
    InMux I__3344 (
            .O(N__19925),
            .I(N__19912));
    InMux I__3343 (
            .O(N__19922),
            .I(N__19907));
    LocalMux I__3342 (
            .O(N__19919),
            .I(N__19903));
    LocalMux I__3341 (
            .O(N__19916),
            .I(N__19900));
    InMux I__3340 (
            .O(N__19915),
            .I(N__19897));
    LocalMux I__3339 (
            .O(N__19912),
            .I(N__19894));
    InMux I__3338 (
            .O(N__19911),
            .I(N__19891));
    InMux I__3337 (
            .O(N__19910),
            .I(N__19888));
    LocalMux I__3336 (
            .O(N__19907),
            .I(N__19885));
    InMux I__3335 (
            .O(N__19906),
            .I(N__19882));
    Span4Mux_h I__3334 (
            .O(N__19903),
            .I(N__19875));
    Span4Mux_v I__3333 (
            .O(N__19900),
            .I(N__19875));
    LocalMux I__3332 (
            .O(N__19897),
            .I(N__19875));
    Span4Mux_h I__3331 (
            .O(N__19894),
            .I(N__19872));
    LocalMux I__3330 (
            .O(N__19891),
            .I(N__19869));
    LocalMux I__3329 (
            .O(N__19888),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv12 I__3328 (
            .O(N__19885),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    LocalMux I__3327 (
            .O(N__19882),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__3326 (
            .O(N__19875),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__3325 (
            .O(N__19872),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    Odrv4 I__3324 (
            .O(N__19869),
            .I(\this_spr_ram.mem_radregZ0Z_11 ));
    InMux I__3323 (
            .O(N__19856),
            .I(N__19853));
    LocalMux I__3322 (
            .O(N__19853),
            .I(\this_ppu.N_797 ));
    InMux I__3321 (
            .O(N__19850),
            .I(N__19847));
    LocalMux I__3320 (
            .O(N__19847),
            .I(M_this_data_tmp_qZ0Z_2));
    InMux I__3319 (
            .O(N__19844),
            .I(N__19841));
    LocalMux I__3318 (
            .O(N__19841),
            .I(N__19838));
    Odrv4 I__3317 (
            .O(N__19838),
            .I(M_this_data_tmp_qZ0Z_21));
    InMux I__3316 (
            .O(N__19835),
            .I(N__19832));
    LocalMux I__3315 (
            .O(N__19832),
            .I(N__19829));
    Span4Mux_v I__3314 (
            .O(N__19829),
            .I(N__19826));
    Span4Mux_v I__3313 (
            .O(N__19826),
            .I(N__19823));
    Span4Mux_v I__3312 (
            .O(N__19823),
            .I(N__19820));
    Span4Mux_v I__3311 (
            .O(N__19820),
            .I(N__19817));
    Span4Mux_h I__3310 (
            .O(N__19817),
            .I(N__19814));
    Odrv4 I__3309 (
            .O(N__19814),
            .I(\this_spr_ram.mem_out_bus7_0 ));
    InMux I__3308 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__3307 (
            .O(N__19808),
            .I(N__19805));
    Span4Mux_h I__3306 (
            .O(N__19805),
            .I(N__19802));
    Span4Mux_h I__3305 (
            .O(N__19802),
            .I(N__19799));
    Span4Mux_h I__3304 (
            .O(N__19799),
            .I(N__19796));
    Odrv4 I__3303 (
            .O(N__19796),
            .I(\this_spr_ram.mem_out_bus3_0 ));
    InMux I__3302 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__3301 (
            .O(N__19790),
            .I(N__19787));
    Span12Mux_v I__3300 (
            .O(N__19787),
            .I(N__19784));
    Span12Mux_h I__3299 (
            .O(N__19784),
            .I(N__19781));
    Odrv12 I__3298 (
            .O(N__19781),
            .I(\this_spr_ram.mem_out_bus4_0 ));
    InMux I__3297 (
            .O(N__19778),
            .I(N__19775));
    LocalMux I__3296 (
            .O(N__19775),
            .I(N__19772));
    Span4Mux_v I__3295 (
            .O(N__19772),
            .I(N__19769));
    Span4Mux_h I__3294 (
            .O(N__19769),
            .I(N__19766));
    Odrv4 I__3293 (
            .O(N__19766),
            .I(\this_spr_ram.mem_out_bus0_0 ));
    InMux I__3292 (
            .O(N__19763),
            .I(N__19760));
    LocalMux I__3291 (
            .O(N__19760),
            .I(N__19757));
    Span4Mux_h I__3290 (
            .O(N__19757),
            .I(N__19754));
    Span4Mux_v I__3289 (
            .O(N__19754),
            .I(N__19751));
    Span4Mux_h I__3288 (
            .O(N__19751),
            .I(N__19748));
    Span4Mux_h I__3287 (
            .O(N__19748),
            .I(N__19745));
    Odrv4 I__3286 (
            .O(N__19745),
            .I(\this_spr_ram.mem_out_bus5_0 ));
    InMux I__3285 (
            .O(N__19742),
            .I(N__19739));
    LocalMux I__3284 (
            .O(N__19739),
            .I(N__19736));
    Span4Mux_v I__3283 (
            .O(N__19736),
            .I(N__19733));
    Span4Mux_h I__3282 (
            .O(N__19733),
            .I(N__19730));
    Odrv4 I__3281 (
            .O(N__19730),
            .I(\this_spr_ram.mem_out_bus1_0 ));
    InMux I__3280 (
            .O(N__19727),
            .I(N__19724));
    LocalMux I__3279 (
            .O(N__19724),
            .I(N__19721));
    Sp12to4 I__3278 (
            .O(N__19721),
            .I(N__19718));
    Span12Mux_v I__3277 (
            .O(N__19718),
            .I(N__19715));
    Span12Mux_h I__3276 (
            .O(N__19715),
            .I(N__19712));
    Odrv12 I__3275 (
            .O(N__19712),
            .I(\this_spr_ram.mem_out_bus6_0 ));
    InMux I__3274 (
            .O(N__19709),
            .I(N__19706));
    LocalMux I__3273 (
            .O(N__19706),
            .I(N__19703));
    Span12Mux_v I__3272 (
            .O(N__19703),
            .I(N__19700));
    Span12Mux_h I__3271 (
            .O(N__19700),
            .I(N__19697));
    Odrv12 I__3270 (
            .O(N__19697),
            .I(\this_spr_ram.mem_out_bus2_0 ));
    CascadeMux I__3269 (
            .O(N__19694),
            .I(N__19689));
    CascadeMux I__3268 (
            .O(N__19693),
            .I(N__19686));
    InMux I__3267 (
            .O(N__19692),
            .I(N__19683));
    InMux I__3266 (
            .O(N__19689),
            .I(N__19679));
    InMux I__3265 (
            .O(N__19686),
            .I(N__19676));
    LocalMux I__3264 (
            .O(N__19683),
            .I(N__19673));
    InMux I__3263 (
            .O(N__19682),
            .I(N__19670));
    LocalMux I__3262 (
            .O(N__19679),
            .I(N__19665));
    LocalMux I__3261 (
            .O(N__19676),
            .I(N__19665));
    Span4Mux_v I__3260 (
            .O(N__19673),
            .I(N__19662));
    LocalMux I__3259 (
            .O(N__19670),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    Odrv12 I__3258 (
            .O(N__19665),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    Odrv4 I__3257 (
            .O(N__19662),
            .I(\this_spr_ram.mem_radregZ0Z_12 ));
    CascadeMux I__3256 (
            .O(N__19655),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ));
    InMux I__3255 (
            .O(N__19652),
            .I(N__19649));
    LocalMux I__3254 (
            .O(N__19649),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ));
    InMux I__3253 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__3252 (
            .O(N__19643),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ));
    InMux I__3251 (
            .O(N__19640),
            .I(N__19637));
    LocalMux I__3250 (
            .O(N__19637),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ));
    InMux I__3249 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__3248 (
            .O(N__19631),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ));
    InMux I__3247 (
            .O(N__19628),
            .I(N__19624));
    InMux I__3246 (
            .O(N__19627),
            .I(N__19621));
    LocalMux I__3245 (
            .O(N__19624),
            .I(N__19618));
    LocalMux I__3244 (
            .O(N__19621),
            .I(N__19615));
    Span4Mux_v I__3243 (
            .O(N__19618),
            .I(N__19612));
    Span4Mux_v I__3242 (
            .O(N__19615),
            .I(N__19609));
    Odrv4 I__3241 (
            .O(N__19612),
            .I(M_this_spr_ram_read_data_0));
    Odrv4 I__3240 (
            .O(N__19609),
            .I(M_this_spr_ram_read_data_0));
    CascadeMux I__3239 (
            .O(N__19604),
            .I(N__19601));
    CascadeBuf I__3238 (
            .O(N__19601),
            .I(N__19598));
    CascadeMux I__3237 (
            .O(N__19598),
            .I(N__19595));
    InMux I__3236 (
            .O(N__19595),
            .I(N__19591));
    CascadeMux I__3235 (
            .O(N__19594),
            .I(N__19588));
    LocalMux I__3234 (
            .O(N__19591),
            .I(N__19584));
    InMux I__3233 (
            .O(N__19588),
            .I(N__19581));
    InMux I__3232 (
            .O(N__19587),
            .I(N__19578));
    Span12Mux_s7_v I__3231 (
            .O(N__19584),
            .I(N__19575));
    LocalMux I__3230 (
            .O(N__19581),
            .I(M_this_oam_address_qZ0Z_3));
    LocalMux I__3229 (
            .O(N__19578),
            .I(M_this_oam_address_qZ0Z_3));
    Odrv12 I__3228 (
            .O(N__19575),
            .I(M_this_oam_address_qZ0Z_3));
    CascadeMux I__3227 (
            .O(N__19568),
            .I(N__19565));
    CascadeBuf I__3226 (
            .O(N__19565),
            .I(N__19562));
    CascadeMux I__3225 (
            .O(N__19562),
            .I(N__19559));
    InMux I__3224 (
            .O(N__19559),
            .I(N__19556));
    LocalMux I__3223 (
            .O(N__19556),
            .I(N__19553));
    Span4Mux_h I__3222 (
            .O(N__19553),
            .I(N__19547));
    InMux I__3221 (
            .O(N__19552),
            .I(N__19542));
    InMux I__3220 (
            .O(N__19551),
            .I(N__19542));
    InMux I__3219 (
            .O(N__19550),
            .I(N__19539));
    Span4Mux_v I__3218 (
            .O(N__19547),
            .I(N__19536));
    LocalMux I__3217 (
            .O(N__19542),
            .I(M_this_oam_address_qZ0Z_2));
    LocalMux I__3216 (
            .O(N__19539),
            .I(M_this_oam_address_qZ0Z_2));
    Odrv4 I__3215 (
            .O(N__19536),
            .I(M_this_oam_address_qZ0Z_2));
    InMux I__3214 (
            .O(N__19529),
            .I(N__19523));
    InMux I__3213 (
            .O(N__19528),
            .I(N__19523));
    LocalMux I__3212 (
            .O(N__19523),
            .I(un1_M_this_oam_address_q_c4));
    CascadeMux I__3211 (
            .O(N__19520),
            .I(N__19517));
    CascadeBuf I__3210 (
            .O(N__19517),
            .I(N__19514));
    CascadeMux I__3209 (
            .O(N__19514),
            .I(N__19511));
    InMux I__3208 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__3207 (
            .O(N__19508),
            .I(N__19505));
    Span4Mux_h I__3206 (
            .O(N__19505),
            .I(N__19500));
    InMux I__3205 (
            .O(N__19504),
            .I(N__19497));
    InMux I__3204 (
            .O(N__19503),
            .I(N__19494));
    Span4Mux_v I__3203 (
            .O(N__19500),
            .I(N__19491));
    LocalMux I__3202 (
            .O(N__19497),
            .I(M_this_oam_address_qZ0Z_5));
    LocalMux I__3201 (
            .O(N__19494),
            .I(M_this_oam_address_qZ0Z_5));
    Odrv4 I__3200 (
            .O(N__19491),
            .I(M_this_oam_address_qZ0Z_5));
    CascadeMux I__3199 (
            .O(N__19484),
            .I(un1_M_this_oam_address_q_c4_cascade_));
    CascadeMux I__3198 (
            .O(N__19481),
            .I(N__19478));
    CascadeBuf I__3197 (
            .O(N__19478),
            .I(N__19475));
    CascadeMux I__3196 (
            .O(N__19475),
            .I(N__19472));
    InMux I__3195 (
            .O(N__19472),
            .I(N__19469));
    LocalMux I__3194 (
            .O(N__19469),
            .I(N__19465));
    CascadeMux I__3193 (
            .O(N__19468),
            .I(N__19462));
    Span4Mux_h I__3192 (
            .O(N__19465),
            .I(N__19457));
    InMux I__3191 (
            .O(N__19462),
            .I(N__19454));
    InMux I__3190 (
            .O(N__19461),
            .I(N__19451));
    InMux I__3189 (
            .O(N__19460),
            .I(N__19448));
    Span4Mux_v I__3188 (
            .O(N__19457),
            .I(N__19445));
    LocalMux I__3187 (
            .O(N__19454),
            .I(M_this_oam_address_qZ0Z_4));
    LocalMux I__3186 (
            .O(N__19451),
            .I(M_this_oam_address_qZ0Z_4));
    LocalMux I__3185 (
            .O(N__19448),
            .I(M_this_oam_address_qZ0Z_4));
    Odrv4 I__3184 (
            .O(N__19445),
            .I(M_this_oam_address_qZ0Z_4));
    InMux I__3183 (
            .O(N__19436),
            .I(N__19430));
    InMux I__3182 (
            .O(N__19435),
            .I(N__19430));
    LocalMux I__3181 (
            .O(N__19430),
            .I(un1_M_this_oam_address_q_c6));
    CEMux I__3180 (
            .O(N__19427),
            .I(N__19423));
    CEMux I__3179 (
            .O(N__19426),
            .I(N__19420));
    LocalMux I__3178 (
            .O(N__19423),
            .I(N__19417));
    LocalMux I__3177 (
            .O(N__19420),
            .I(N__19414));
    Odrv4 I__3176 (
            .O(N__19417),
            .I(N_1240_0));
    Odrv12 I__3175 (
            .O(N__19414),
            .I(N_1240_0));
    CascadeMux I__3174 (
            .O(N__19409),
            .I(M_this_oam_ram_write_data_0_sqmuxa_cascade_));
    InMux I__3173 (
            .O(N__19406),
            .I(N__19403));
    LocalMux I__3172 (
            .O(N__19403),
            .I(N__19400));
    Span4Mux_s2_v I__3171 (
            .O(N__19400),
            .I(N__19397));
    Span4Mux_h I__3170 (
            .O(N__19397),
            .I(N__19394));
    Odrv4 I__3169 (
            .O(N__19394),
            .I(M_this_oam_ram_write_data_26));
    CEMux I__3168 (
            .O(N__19391),
            .I(N__19387));
    CEMux I__3167 (
            .O(N__19390),
            .I(N__19366));
    LocalMux I__3166 (
            .O(N__19387),
            .I(N__19359));
    InMux I__3165 (
            .O(N__19386),
            .I(N__19352));
    InMux I__3164 (
            .O(N__19385),
            .I(N__19352));
    InMux I__3163 (
            .O(N__19384),
            .I(N__19352));
    InMux I__3162 (
            .O(N__19383),
            .I(N__19341));
    InMux I__3161 (
            .O(N__19382),
            .I(N__19341));
    InMux I__3160 (
            .O(N__19381),
            .I(N__19341));
    InMux I__3159 (
            .O(N__19380),
            .I(N__19341));
    InMux I__3158 (
            .O(N__19379),
            .I(N__19341));
    InMux I__3157 (
            .O(N__19378),
            .I(N__19338));
    InMux I__3156 (
            .O(N__19377),
            .I(N__19329));
    InMux I__3155 (
            .O(N__19376),
            .I(N__19329));
    InMux I__3154 (
            .O(N__19375),
            .I(N__19329));
    InMux I__3153 (
            .O(N__19374),
            .I(N__19329));
    InMux I__3152 (
            .O(N__19373),
            .I(N__19316));
    InMux I__3151 (
            .O(N__19372),
            .I(N__19316));
    InMux I__3150 (
            .O(N__19371),
            .I(N__19316));
    InMux I__3149 (
            .O(N__19370),
            .I(N__19316));
    InMux I__3148 (
            .O(N__19369),
            .I(N__19316));
    LocalMux I__3147 (
            .O(N__19366),
            .I(N__19313));
    InMux I__3146 (
            .O(N__19365),
            .I(N__19310));
    InMux I__3145 (
            .O(N__19364),
            .I(N__19307));
    InMux I__3144 (
            .O(N__19363),
            .I(N__19302));
    InMux I__3143 (
            .O(N__19362),
            .I(N__19302));
    Span4Mux_h I__3142 (
            .O(N__19359),
            .I(N__19291));
    LocalMux I__3141 (
            .O(N__19352),
            .I(N__19291));
    LocalMux I__3140 (
            .O(N__19341),
            .I(N__19284));
    LocalMux I__3139 (
            .O(N__19338),
            .I(N__19284));
    LocalMux I__3138 (
            .O(N__19329),
            .I(N__19284));
    InMux I__3137 (
            .O(N__19328),
            .I(N__19279));
    InMux I__3136 (
            .O(N__19327),
            .I(N__19279));
    LocalMux I__3135 (
            .O(N__19316),
            .I(N__19276));
    Span4Mux_h I__3134 (
            .O(N__19313),
            .I(N__19267));
    LocalMux I__3133 (
            .O(N__19310),
            .I(N__19267));
    LocalMux I__3132 (
            .O(N__19307),
            .I(N__19267));
    LocalMux I__3131 (
            .O(N__19302),
            .I(N__19267));
    InMux I__3130 (
            .O(N__19301),
            .I(N__19253));
    InMux I__3129 (
            .O(N__19300),
            .I(N__19253));
    InMux I__3128 (
            .O(N__19299),
            .I(N__19253));
    InMux I__3127 (
            .O(N__19298),
            .I(N__19253));
    InMux I__3126 (
            .O(N__19297),
            .I(N__19253));
    InMux I__3125 (
            .O(N__19296),
            .I(N__19253));
    Span4Mux_s2_v I__3124 (
            .O(N__19291),
            .I(N__19250));
    Span4Mux_v I__3123 (
            .O(N__19284),
            .I(N__19241));
    LocalMux I__3122 (
            .O(N__19279),
            .I(N__19241));
    Span4Mux_h I__3121 (
            .O(N__19276),
            .I(N__19241));
    Span4Mux_v I__3120 (
            .O(N__19267),
            .I(N__19241));
    InMux I__3119 (
            .O(N__19266),
            .I(N__19238));
    LocalMux I__3118 (
            .O(N__19253),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__3117 (
            .O(N__19250),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    Odrv4 I__3116 (
            .O(N__19241),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    LocalMux I__3115 (
            .O(N__19238),
            .I(M_this_oam_ram_write_data_0_sqmuxa));
    InMux I__3114 (
            .O(N__19229),
            .I(N__19226));
    LocalMux I__3113 (
            .O(N__19226),
            .I(N__19223));
    Span4Mux_s3_v I__3112 (
            .O(N__19223),
            .I(N__19220));
    Span4Mux_h I__3111 (
            .O(N__19220),
            .I(N__19217));
    Odrv4 I__3110 (
            .O(N__19217),
            .I(M_this_oam_ram_write_data_0));
    InMux I__3109 (
            .O(N__19214),
            .I(N__19211));
    LocalMux I__3108 (
            .O(N__19211),
            .I(M_this_data_tmp_qZ0Z_0));
    InMux I__3107 (
            .O(N__19208),
            .I(N__19205));
    LocalMux I__3106 (
            .O(N__19205),
            .I(M_this_data_tmp_qZ0Z_4));
    InMux I__3105 (
            .O(N__19202),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_6 ));
    InMux I__3104 (
            .O(N__19199),
            .I(N__19196));
    LocalMux I__3103 (
            .O(N__19196),
            .I(\this_ppu.M_state_q_RNISP3R6_1Z0Z_10 ));
    InMux I__3102 (
            .O(N__19193),
            .I(N__19190));
    LocalMux I__3101 (
            .O(N__19190),
            .I(N__19187));
    Span12Mux_h I__3100 (
            .O(N__19187),
            .I(N__19184));
    Odrv12 I__3099 (
            .O(N__19184),
            .I(M_this_oam_ram_read_data_11));
    InMux I__3098 (
            .O(N__19181),
            .I(N__19178));
    LocalMux I__3097 (
            .O(N__19178),
            .I(N__19175));
    Span4Mux_v I__3096 (
            .O(N__19175),
            .I(N__19172));
    Span4Mux_h I__3095 (
            .O(N__19172),
            .I(N__19169));
    Odrv4 I__3094 (
            .O(N__19169),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_11 ));
    InMux I__3093 (
            .O(N__19166),
            .I(N__19163));
    LocalMux I__3092 (
            .O(N__19163),
            .I(\this_ppu.M_state_q_RNISP3R6Z0Z_10 ));
    InMux I__3091 (
            .O(N__19160),
            .I(N__19152));
    InMux I__3090 (
            .O(N__19159),
            .I(N__19149));
    InMux I__3089 (
            .O(N__19158),
            .I(N__19140));
    InMux I__3088 (
            .O(N__19157),
            .I(N__19140));
    InMux I__3087 (
            .O(N__19156),
            .I(N__19140));
    InMux I__3086 (
            .O(N__19155),
            .I(N__19140));
    LocalMux I__3085 (
            .O(N__19152),
            .I(\this_ppu.N_806 ));
    LocalMux I__3084 (
            .O(N__19149),
            .I(\this_ppu.N_806 ));
    LocalMux I__3083 (
            .O(N__19140),
            .I(\this_ppu.N_806 ));
    InMux I__3082 (
            .O(N__19133),
            .I(N__19130));
    LocalMux I__3081 (
            .O(N__19130),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1 ));
    InMux I__3080 (
            .O(N__19127),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_0 ));
    InMux I__3079 (
            .O(N__19124),
            .I(N__19121));
    LocalMux I__3078 (
            .O(N__19121),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2 ));
    InMux I__3077 (
            .O(N__19118),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_1 ));
    InMux I__3076 (
            .O(N__19115),
            .I(N__19111));
    InMux I__3075 (
            .O(N__19114),
            .I(N__19108));
    LocalMux I__3074 (
            .O(N__19111),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_3 ));
    LocalMux I__3073 (
            .O(N__19108),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_3 ));
    InMux I__3072 (
            .O(N__19103),
            .I(N__19100));
    LocalMux I__3071 (
            .O(N__19100),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3 ));
    InMux I__3070 (
            .O(N__19097),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_2 ));
    CascadeMux I__3069 (
            .O(N__19094),
            .I(N__19091));
    InMux I__3068 (
            .O(N__19091),
            .I(N__19087));
    InMux I__3067 (
            .O(N__19090),
            .I(N__19084));
    LocalMux I__3066 (
            .O(N__19087),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_4 ));
    LocalMux I__3065 (
            .O(N__19084),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_4 ));
    InMux I__3064 (
            .O(N__19079),
            .I(N__19076));
    LocalMux I__3063 (
            .O(N__19076),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4 ));
    InMux I__3062 (
            .O(N__19073),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_3 ));
    CascadeMux I__3061 (
            .O(N__19070),
            .I(N__19067));
    InMux I__3060 (
            .O(N__19067),
            .I(N__19063));
    InMux I__3059 (
            .O(N__19066),
            .I(N__19060));
    LocalMux I__3058 (
            .O(N__19063),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_5 ));
    LocalMux I__3057 (
            .O(N__19060),
            .I(\this_ppu.M_pixel_cnt_qZ1Z_5 ));
    InMux I__3056 (
            .O(N__19055),
            .I(N__19052));
    LocalMux I__3055 (
            .O(N__19052),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5 ));
    InMux I__3054 (
            .O(N__19049),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_4 ));
    CascadeMux I__3053 (
            .O(N__19046),
            .I(N__19043));
    InMux I__3052 (
            .O(N__19043),
            .I(N__19039));
    CascadeMux I__3051 (
            .O(N__19042),
            .I(N__19036));
    LocalMux I__3050 (
            .O(N__19039),
            .I(N__19033));
    InMux I__3049 (
            .O(N__19036),
            .I(N__19030));
    Odrv4 I__3048 (
            .O(N__19033),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_6 ));
    LocalMux I__3047 (
            .O(N__19030),
            .I(\this_ppu.M_pixel_cnt_qZ0Z_6 ));
    InMux I__3046 (
            .O(N__19025),
            .I(N__19022));
    LocalMux I__3045 (
            .O(N__19022),
            .I(N__19019));
    Span4Mux_h I__3044 (
            .O(N__19019),
            .I(N__19016));
    Odrv4 I__3043 (
            .O(N__19016),
            .I(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6 ));
    InMux I__3042 (
            .O(N__19013),
            .I(\this_ppu.un1_M_pixel_cnt_q_1_cry_5 ));
    CascadeMux I__3041 (
            .O(N__19010),
            .I(\this_ppu.m9_0_a2_5_cascade_ ));
    InMux I__3040 (
            .O(N__19007),
            .I(N__19004));
    LocalMux I__3039 (
            .O(N__19004),
            .I(\this_vga_signals.i22_mux ));
    InMux I__3038 (
            .O(N__19001),
            .I(N__18997));
    InMux I__3037 (
            .O(N__19000),
            .I(N__18993));
    LocalMux I__3036 (
            .O(N__18997),
            .I(N__18990));
    InMux I__3035 (
            .O(N__18996),
            .I(N__18987));
    LocalMux I__3034 (
            .O(N__18993),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    Odrv4 I__3033 (
            .O(N__18990),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    LocalMux I__3032 (
            .O(N__18987),
            .I(\this_vga_signals.M_lcounter_qZ0Z_1 ));
    InMux I__3031 (
            .O(N__18980),
            .I(N__18971));
    InMux I__3030 (
            .O(N__18979),
            .I(N__18971));
    InMux I__3029 (
            .O(N__18978),
            .I(N__18971));
    LocalMux I__3028 (
            .O(N__18971),
            .I(\this_vga_signals.M_lcounter_qZ0Z_0 ));
    InMux I__3027 (
            .O(N__18968),
            .I(N__18965));
    LocalMux I__3026 (
            .O(N__18965),
            .I(\this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2 ));
    CascadeMux I__3025 (
            .O(N__18962),
            .I(\this_ppu.N_814_cascade_ ));
    CascadeMux I__3024 (
            .O(N__18959),
            .I(\this_ppu.N_806_cascade_ ));
    InMux I__3023 (
            .O(N__18956),
            .I(N__18950));
    InMux I__3022 (
            .O(N__18955),
            .I(N__18950));
    LocalMux I__3021 (
            .O(N__18950),
            .I(\this_ppu.un1_M_oam_curr_q_1_c5 ));
    CascadeMux I__3020 (
            .O(N__18947),
            .I(N__18944));
    CascadeBuf I__3019 (
            .O(N__18944),
            .I(N__18941));
    CascadeMux I__3018 (
            .O(N__18941),
            .I(N__18938));
    InMux I__3017 (
            .O(N__18938),
            .I(N__18935));
    LocalMux I__3016 (
            .O(N__18935),
            .I(N__18932));
    Span4Mux_h I__3015 (
            .O(N__18932),
            .I(N__18929));
    Span4Mux_v I__3014 (
            .O(N__18929),
            .I(N__18923));
    CascadeMux I__3013 (
            .O(N__18928),
            .I(N__18920));
    InMux I__3012 (
            .O(N__18927),
            .I(N__18917));
    CascadeMux I__3011 (
            .O(N__18926),
            .I(N__18914));
    Span4Mux_v I__3010 (
            .O(N__18923),
            .I(N__18911));
    InMux I__3009 (
            .O(N__18920),
            .I(N__18908));
    LocalMux I__3008 (
            .O(N__18917),
            .I(N__18905));
    InMux I__3007 (
            .O(N__18914),
            .I(N__18902));
    Span4Mux_v I__3006 (
            .O(N__18911),
            .I(N__18899));
    LocalMux I__3005 (
            .O(N__18908),
            .I(M_this_ppu_oam_addr_5));
    Odrv4 I__3004 (
            .O(N__18905),
            .I(M_this_ppu_oam_addr_5));
    LocalMux I__3003 (
            .O(N__18902),
            .I(M_this_ppu_oam_addr_5));
    Odrv4 I__3002 (
            .O(N__18899),
            .I(M_this_ppu_oam_addr_5));
    InMux I__3001 (
            .O(N__18890),
            .I(N__18882));
    InMux I__3000 (
            .O(N__18889),
            .I(N__18877));
    InMux I__2999 (
            .O(N__18888),
            .I(N__18877));
    InMux I__2998 (
            .O(N__18887),
            .I(N__18874));
    InMux I__2997 (
            .O(N__18886),
            .I(N__18869));
    InMux I__2996 (
            .O(N__18885),
            .I(N__18869));
    LocalMux I__2995 (
            .O(N__18882),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    LocalMux I__2994 (
            .O(N__18877),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    LocalMux I__2993 (
            .O(N__18874),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    LocalMux I__2992 (
            .O(N__18869),
            .I(\this_ppu.M_oam_curr_qc_0_1 ));
    InMux I__2991 (
            .O(N__18860),
            .I(N__18856));
    InMux I__2990 (
            .O(N__18859),
            .I(N__18853));
    LocalMux I__2989 (
            .O(N__18856),
            .I(N__18850));
    LocalMux I__2988 (
            .O(N__18853),
            .I(\this_ppu.M_oam_curr_qZ0Z_6 ));
    Odrv4 I__2987 (
            .O(N__18850),
            .I(\this_ppu.M_oam_curr_qZ0Z_6 ));
    InMux I__2986 (
            .O(N__18845),
            .I(N__18842));
    LocalMux I__2985 (
            .O(N__18842),
            .I(N__18838));
    CascadeMux I__2984 (
            .O(N__18841),
            .I(N__18835));
    Span4Mux_h I__2983 (
            .O(N__18838),
            .I(N__18832));
    InMux I__2982 (
            .O(N__18835),
            .I(N__18828));
    Span4Mux_v I__2981 (
            .O(N__18832),
            .I(N__18825));
    InMux I__2980 (
            .O(N__18831),
            .I(N__18822));
    LocalMux I__2979 (
            .O(N__18828),
            .I(N__18819));
    Odrv4 I__2978 (
            .O(N__18825),
            .I(M_this_status_flags_qZ0Z_0));
    LocalMux I__2977 (
            .O(N__18822),
            .I(M_this_status_flags_qZ0Z_0));
    Odrv12 I__2976 (
            .O(N__18819),
            .I(M_this_status_flags_qZ0Z_0));
    InMux I__2975 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__2974 (
            .O(N__18809),
            .I(N__18806));
    Span4Mux_h I__2973 (
            .O(N__18806),
            .I(N__18803));
    Odrv4 I__2972 (
            .O(N__18803),
            .I(\this_ppu.oam_cache.mem_15 ));
    InMux I__2971 (
            .O(N__18800),
            .I(N__18791));
    InMux I__2970 (
            .O(N__18799),
            .I(N__18791));
    InMux I__2969 (
            .O(N__18798),
            .I(N__18791));
    LocalMux I__2968 (
            .O(N__18791),
            .I(N__18788));
    Span4Mux_h I__2967 (
            .O(N__18788),
            .I(N__18784));
    InMux I__2966 (
            .O(N__18787),
            .I(N__18781));
    Odrv4 I__2965 (
            .O(N__18784),
            .I(\this_ppu.N_784_0 ));
    LocalMux I__2964 (
            .O(N__18781),
            .I(\this_ppu.N_784_0 ));
    CascadeMux I__2963 (
            .O(N__18776),
            .I(\this_vga_signals.N_859_cascade_ ));
    InMux I__2962 (
            .O(N__18773),
            .I(N__18770));
    LocalMux I__2961 (
            .O(N__18770),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_13 ));
    InMux I__2960 (
            .O(N__18767),
            .I(N__18764));
    LocalMux I__2959 (
            .O(N__18764),
            .I(\this_spr_ram.mem_mem_3_1_RNISI5GZ0 ));
    CascadeMux I__2958 (
            .O(N__18761),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ));
    InMux I__2957 (
            .O(N__18758),
            .I(N__18755));
    LocalMux I__2956 (
            .O(N__18755),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ));
    CascadeMux I__2955 (
            .O(N__18752),
            .I(N__18749));
    InMux I__2954 (
            .O(N__18749),
            .I(N__18743));
    InMux I__2953 (
            .O(N__18748),
            .I(N__18740));
    InMux I__2952 (
            .O(N__18747),
            .I(N__18737));
    InMux I__2951 (
            .O(N__18746),
            .I(N__18734));
    LocalMux I__2950 (
            .O(N__18743),
            .I(N__18731));
    LocalMux I__2949 (
            .O(N__18740),
            .I(N__18726));
    LocalMux I__2948 (
            .O(N__18737),
            .I(N__18726));
    LocalMux I__2947 (
            .O(N__18734),
            .I(N__18723));
    Span4Mux_h I__2946 (
            .O(N__18731),
            .I(N__18718));
    Span4Mux_v I__2945 (
            .O(N__18726),
            .I(N__18718));
    Span4Mux_v I__2944 (
            .O(N__18723),
            .I(N__18713));
    Span4Mux_v I__2943 (
            .O(N__18718),
            .I(N__18713));
    Odrv4 I__2942 (
            .O(N__18713),
            .I(this_ppu_N_247));
    InMux I__2941 (
            .O(N__18710),
            .I(N__18707));
    LocalMux I__2940 (
            .O(N__18707),
            .I(N__18703));
    InMux I__2939 (
            .O(N__18706),
            .I(N__18700));
    Odrv4 I__2938 (
            .O(N__18703),
            .I(\this_vga_signals.N_22_0 ));
    LocalMux I__2937 (
            .O(N__18700),
            .I(\this_vga_signals.N_22_0 ));
    CascadeMux I__2936 (
            .O(N__18695),
            .I(M_this_spr_ram_read_data_2_cascade_));
    InMux I__2935 (
            .O(N__18692),
            .I(N__18689));
    LocalMux I__2934 (
            .O(N__18689),
            .I(N__18686));
    Span4Mux_h I__2933 (
            .O(N__18686),
            .I(N__18683));
    Odrv4 I__2932 (
            .O(N__18683),
            .I(N_28_0_i));
    CascadeMux I__2931 (
            .O(N__18680),
            .I(N__18677));
    CascadeBuf I__2930 (
            .O(N__18677),
            .I(N__18674));
    CascadeMux I__2929 (
            .O(N__18674),
            .I(N__18671));
    InMux I__2928 (
            .O(N__18671),
            .I(N__18667));
    InMux I__2927 (
            .O(N__18670),
            .I(N__18663));
    LocalMux I__2926 (
            .O(N__18667),
            .I(N__18660));
    InMux I__2925 (
            .O(N__18666),
            .I(N__18657));
    LocalMux I__2924 (
            .O(N__18663),
            .I(N__18654));
    Span4Mux_h I__2923 (
            .O(N__18660),
            .I(N__18651));
    LocalMux I__2922 (
            .O(N__18657),
            .I(N__18647));
    Span4Mux_h I__2921 (
            .O(N__18654),
            .I(N__18643));
    Sp12to4 I__2920 (
            .O(N__18651),
            .I(N__18640));
    InMux I__2919 (
            .O(N__18650),
            .I(N__18637));
    Span4Mux_h I__2918 (
            .O(N__18647),
            .I(N__18634));
    InMux I__2917 (
            .O(N__18646),
            .I(N__18631));
    Sp12to4 I__2916 (
            .O(N__18643),
            .I(N__18626));
    Span12Mux_s7_v I__2915 (
            .O(N__18640),
            .I(N__18626));
    LocalMux I__2914 (
            .O(N__18637),
            .I(M_this_ppu_oam_addr_4));
    Odrv4 I__2913 (
            .O(N__18634),
            .I(M_this_ppu_oam_addr_4));
    LocalMux I__2912 (
            .O(N__18631),
            .I(M_this_ppu_oam_addr_4));
    Odrv12 I__2911 (
            .O(N__18626),
            .I(M_this_ppu_oam_addr_4));
    InMux I__2910 (
            .O(N__18617),
            .I(N__18614));
    LocalMux I__2909 (
            .O(N__18614),
            .I(M_this_spr_ram_read_data_2));
    InMux I__2908 (
            .O(N__18611),
            .I(N__18607));
    InMux I__2907 (
            .O(N__18610),
            .I(N__18604));
    LocalMux I__2906 (
            .O(N__18607),
            .I(N__18599));
    LocalMux I__2905 (
            .O(N__18604),
            .I(N__18599));
    Odrv12 I__2904 (
            .O(N__18599),
            .I(M_this_spr_ram_read_data_1));
    CascadeMux I__2903 (
            .O(N__18596),
            .I(N__18593));
    InMux I__2902 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__2901 (
            .O(N__18590),
            .I(N__18587));
    Span4Mux_h I__2900 (
            .O(N__18587),
            .I(N__18584));
    Odrv4 I__2899 (
            .O(N__18584),
            .I(M_this_spr_ram_read_data_3));
    CascadeMux I__2898 (
            .O(N__18581),
            .I(\this_ppu.M_oam_curr_dZ0Z25_cascade_ ));
    InMux I__2897 (
            .O(N__18578),
            .I(N__18575));
    LocalMux I__2896 (
            .O(N__18575),
            .I(N__18572));
    Span4Mux_h I__2895 (
            .O(N__18572),
            .I(N__18567));
    InMux I__2894 (
            .O(N__18571),
            .I(N__18564));
    InMux I__2893 (
            .O(N__18570),
            .I(N__18561));
    Span4Mux_v I__2892 (
            .O(N__18567),
            .I(N__18558));
    LocalMux I__2891 (
            .O(N__18564),
            .I(\this_ppu.N_834_0 ));
    LocalMux I__2890 (
            .O(N__18561),
            .I(\this_ppu.N_834_0 ));
    Odrv4 I__2889 (
            .O(N__18558),
            .I(\this_ppu.N_834_0 ));
    CascadeMux I__2888 (
            .O(N__18551),
            .I(N__18548));
    CascadeBuf I__2887 (
            .O(N__18548),
            .I(N__18545));
    CascadeMux I__2886 (
            .O(N__18545),
            .I(N__18541));
    InMux I__2885 (
            .O(N__18544),
            .I(N__18537));
    InMux I__2884 (
            .O(N__18541),
            .I(N__18534));
    InMux I__2883 (
            .O(N__18540),
            .I(N__18530));
    LocalMux I__2882 (
            .O(N__18537),
            .I(N__18527));
    LocalMux I__2881 (
            .O(N__18534),
            .I(N__18524));
    CascadeMux I__2880 (
            .O(N__18533),
            .I(N__18521));
    LocalMux I__2879 (
            .O(N__18530),
            .I(N__18518));
    Span4Mux_v I__2878 (
            .O(N__18527),
            .I(N__18514));
    Span12Mux_s10_h I__2877 (
            .O(N__18524),
            .I(N__18510));
    InMux I__2876 (
            .O(N__18521),
            .I(N__18507));
    Span4Mux_v I__2875 (
            .O(N__18518),
            .I(N__18504));
    InMux I__2874 (
            .O(N__18517),
            .I(N__18501));
    Span4Mux_h I__2873 (
            .O(N__18514),
            .I(N__18498));
    InMux I__2872 (
            .O(N__18513),
            .I(N__18495));
    Span12Mux_v I__2871 (
            .O(N__18510),
            .I(N__18492));
    LocalMux I__2870 (
            .O(N__18507),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__2869 (
            .O(N__18504),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__2868 (
            .O(N__18501),
            .I(M_this_ppu_oam_addr_0));
    Odrv4 I__2867 (
            .O(N__18498),
            .I(M_this_ppu_oam_addr_0));
    LocalMux I__2866 (
            .O(N__18495),
            .I(M_this_ppu_oam_addr_0));
    Odrv12 I__2865 (
            .O(N__18492),
            .I(M_this_ppu_oam_addr_0));
    CascadeMux I__2864 (
            .O(N__18479),
            .I(\this_ppu.N_834_0_cascade_ ));
    InMux I__2863 (
            .O(N__18476),
            .I(N__18472));
    InMux I__2862 (
            .O(N__18475),
            .I(N__18469));
    LocalMux I__2861 (
            .O(N__18472),
            .I(N__18463));
    LocalMux I__2860 (
            .O(N__18469),
            .I(N__18463));
    InMux I__2859 (
            .O(N__18468),
            .I(N__18460));
    Span4Mux_h I__2858 (
            .O(N__18463),
            .I(N__18457));
    LocalMux I__2857 (
            .O(N__18460),
            .I(\this_ppu.un1_M_state_q_7_i_0_0 ));
    Odrv4 I__2856 (
            .O(N__18457),
            .I(\this_ppu.un1_M_state_q_7_i_0_0 ));
    InMux I__2855 (
            .O(N__18452),
            .I(N__18446));
    InMux I__2854 (
            .O(N__18451),
            .I(N__18446));
    LocalMux I__2853 (
            .O(N__18446),
            .I(N__18441));
    InMux I__2852 (
            .O(N__18445),
            .I(N__18438));
    InMux I__2851 (
            .O(N__18444),
            .I(N__18435));
    Span4Mux_v I__2850 (
            .O(N__18441),
            .I(N__18432));
    LocalMux I__2849 (
            .O(N__18438),
            .I(\this_ppu.un1_M_oam_curr_q_1_c1 ));
    LocalMux I__2848 (
            .O(N__18435),
            .I(\this_ppu.un1_M_oam_curr_q_1_c1 ));
    Odrv4 I__2847 (
            .O(N__18432),
            .I(\this_ppu.un1_M_oam_curr_q_1_c1 ));
    CascadeMux I__2846 (
            .O(N__18425),
            .I(N__18422));
    CascadeBuf I__2845 (
            .O(N__18422),
            .I(N__18419));
    CascadeMux I__2844 (
            .O(N__18419),
            .I(N__18416));
    InMux I__2843 (
            .O(N__18416),
            .I(N__18413));
    LocalMux I__2842 (
            .O(N__18413),
            .I(N__18410));
    Span4Mux_v I__2841 (
            .O(N__18410),
            .I(N__18404));
    InMux I__2840 (
            .O(N__18409),
            .I(N__18399));
    InMux I__2839 (
            .O(N__18408),
            .I(N__18399));
    InMux I__2838 (
            .O(N__18407),
            .I(N__18396));
    Sp12to4 I__2837 (
            .O(N__18404),
            .I(N__18393));
    LocalMux I__2836 (
            .O(N__18399),
            .I(N__18389));
    LocalMux I__2835 (
            .O(N__18396),
            .I(N__18381));
    Span12Mux_s6_h I__2834 (
            .O(N__18393),
            .I(N__18381));
    InMux I__2833 (
            .O(N__18392),
            .I(N__18378));
    Span4Mux_v I__2832 (
            .O(N__18389),
            .I(N__18375));
    InMux I__2831 (
            .O(N__18388),
            .I(N__18370));
    InMux I__2830 (
            .O(N__18387),
            .I(N__18370));
    InMux I__2829 (
            .O(N__18386),
            .I(N__18367));
    Span12Mux_v I__2828 (
            .O(N__18381),
            .I(N__18364));
    LocalMux I__2827 (
            .O(N__18378),
            .I(M_this_ppu_oam_addr_1));
    Odrv4 I__2826 (
            .O(N__18375),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__2825 (
            .O(N__18370),
            .I(M_this_ppu_oam_addr_1));
    LocalMux I__2824 (
            .O(N__18367),
            .I(M_this_ppu_oam_addr_1));
    Odrv12 I__2823 (
            .O(N__18364),
            .I(M_this_ppu_oam_addr_1));
    CascadeMux I__2822 (
            .O(N__18353),
            .I(\this_ppu.un1_M_oam_curr_q_1_c1_cascade_ ));
    CascadeMux I__2821 (
            .O(N__18350),
            .I(N__18346));
    CascadeMux I__2820 (
            .O(N__18349),
            .I(N__18343));
    InMux I__2819 (
            .O(N__18346),
            .I(N__18340));
    CascadeBuf I__2818 (
            .O(N__18343),
            .I(N__18336));
    LocalMux I__2817 (
            .O(N__18340),
            .I(N__18333));
    InMux I__2816 (
            .O(N__18339),
            .I(N__18330));
    CascadeMux I__2815 (
            .O(N__18336),
            .I(N__18327));
    Span4Mux_v I__2814 (
            .O(N__18333),
            .I(N__18324));
    LocalMux I__2813 (
            .O(N__18330),
            .I(N__18321));
    InMux I__2812 (
            .O(N__18327),
            .I(N__18318));
    Sp12to4 I__2811 (
            .O(N__18324),
            .I(N__18314));
    Span4Mux_h I__2810 (
            .O(N__18321),
            .I(N__18311));
    LocalMux I__2809 (
            .O(N__18318),
            .I(N__18308));
    CascadeMux I__2808 (
            .O(N__18317),
            .I(N__18305));
    Span12Mux_h I__2807 (
            .O(N__18314),
            .I(N__18296));
    Sp12to4 I__2806 (
            .O(N__18311),
            .I(N__18296));
    Span12Mux_s10_h I__2805 (
            .O(N__18308),
            .I(N__18296));
    InMux I__2804 (
            .O(N__18305),
            .I(N__18293));
    InMux I__2803 (
            .O(N__18304),
            .I(N__18290));
    InMux I__2802 (
            .O(N__18303),
            .I(N__18287));
    Span12Mux_v I__2801 (
            .O(N__18296),
            .I(N__18284));
    LocalMux I__2800 (
            .O(N__18293),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__2799 (
            .O(N__18290),
            .I(M_this_ppu_oam_addr_2));
    LocalMux I__2798 (
            .O(N__18287),
            .I(M_this_ppu_oam_addr_2));
    Odrv12 I__2797 (
            .O(N__18284),
            .I(M_this_ppu_oam_addr_2));
    InMux I__2796 (
            .O(N__18275),
            .I(N__18268));
    InMux I__2795 (
            .O(N__18274),
            .I(N__18268));
    InMux I__2794 (
            .O(N__18273),
            .I(N__18265));
    LocalMux I__2793 (
            .O(N__18268),
            .I(\this_ppu.un1_M_oam_curr_q_1_c3 ));
    LocalMux I__2792 (
            .O(N__18265),
            .I(\this_ppu.un1_M_oam_curr_q_1_c3 ));
    CascadeMux I__2791 (
            .O(N__18260),
            .I(N__18257));
    CascadeBuf I__2790 (
            .O(N__18257),
            .I(N__18254));
    CascadeMux I__2789 (
            .O(N__18254),
            .I(N__18251));
    InMux I__2788 (
            .O(N__18251),
            .I(N__18248));
    LocalMux I__2787 (
            .O(N__18248),
            .I(N__18244));
    InMux I__2786 (
            .O(N__18247),
            .I(N__18241));
    Span4Mux_v I__2785 (
            .O(N__18244),
            .I(N__18237));
    LocalMux I__2784 (
            .O(N__18241),
            .I(N__18233));
    InMux I__2783 (
            .O(N__18240),
            .I(N__18230));
    Span4Mux_v I__2782 (
            .O(N__18237),
            .I(N__18227));
    CascadeMux I__2781 (
            .O(N__18236),
            .I(N__18224));
    Span4Mux_h I__2780 (
            .O(N__18233),
            .I(N__18218));
    LocalMux I__2779 (
            .O(N__18230),
            .I(N__18213));
    Span4Mux_v I__2778 (
            .O(N__18227),
            .I(N__18213));
    InMux I__2777 (
            .O(N__18224),
            .I(N__18208));
    InMux I__2776 (
            .O(N__18223),
            .I(N__18208));
    InMux I__2775 (
            .O(N__18222),
            .I(N__18203));
    InMux I__2774 (
            .O(N__18221),
            .I(N__18203));
    Span4Mux_v I__2773 (
            .O(N__18218),
            .I(N__18200));
    Span4Mux_v I__2772 (
            .O(N__18213),
            .I(N__18197));
    LocalMux I__2771 (
            .O(N__18208),
            .I(M_this_ppu_oam_addr_3));
    LocalMux I__2770 (
            .O(N__18203),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__2769 (
            .O(N__18200),
            .I(M_this_ppu_oam_addr_3));
    Odrv4 I__2768 (
            .O(N__18197),
            .I(M_this_ppu_oam_addr_3));
    CascadeMux I__2767 (
            .O(N__18188),
            .I(\this_ppu.un1_M_oam_curr_q_1_c3_cascade_ ));
    CascadeMux I__2766 (
            .O(N__18185),
            .I(N__18182));
    CascadeBuf I__2765 (
            .O(N__18182),
            .I(N__18179));
    CascadeMux I__2764 (
            .O(N__18179),
            .I(N__18176));
    InMux I__2763 (
            .O(N__18176),
            .I(N__18173));
    LocalMux I__2762 (
            .O(N__18173),
            .I(N__18170));
    Span4Mux_v I__2761 (
            .O(N__18170),
            .I(N__18167));
    Span4Mux_h I__2760 (
            .O(N__18167),
            .I(N__18164));
    Odrv4 I__2759 (
            .O(N__18164),
            .I(\this_ppu.N_778_0 ));
    InMux I__2758 (
            .O(N__18161),
            .I(N__18158));
    LocalMux I__2757 (
            .O(N__18158),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_14 ));
    InMux I__2756 (
            .O(N__18155),
            .I(N__18152));
    LocalMux I__2755 (
            .O(N__18152),
            .I(N__18149));
    Span4Mux_v I__2754 (
            .O(N__18149),
            .I(N__18146));
    Span4Mux_h I__2753 (
            .O(N__18146),
            .I(N__18143));
    Sp12to4 I__2752 (
            .O(N__18143),
            .I(N__18140));
    Odrv12 I__2751 (
            .O(N__18140),
            .I(\this_spr_ram.mem_out_bus4_2 ));
    InMux I__2750 (
            .O(N__18137),
            .I(N__18134));
    LocalMux I__2749 (
            .O(N__18134),
            .I(N__18131));
    Span12Mux_v I__2748 (
            .O(N__18131),
            .I(N__18128));
    Odrv12 I__2747 (
            .O(N__18128),
            .I(\this_spr_ram.mem_out_bus0_2 ));
    InMux I__2746 (
            .O(N__18125),
            .I(N__18122));
    LocalMux I__2745 (
            .O(N__18122),
            .I(N__18119));
    Span4Mux_h I__2744 (
            .O(N__18119),
            .I(N__18116));
    Odrv4 I__2743 (
            .O(N__18116),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_6 ));
    CascadeMux I__2742 (
            .O(N__18113),
            .I(\this_ppu.M_state_q_inv_1_cascade_ ));
    InMux I__2741 (
            .O(N__18110),
            .I(N__18107));
    LocalMux I__2740 (
            .O(N__18107),
            .I(N__18104));
    Span4Mux_v I__2739 (
            .O(N__18104),
            .I(N__18101));
    Sp12to4 I__2738 (
            .O(N__18101),
            .I(N__18098));
    Span12Mux_h I__2737 (
            .O(N__18098),
            .I(N__18095));
    Span12Mux_v I__2736 (
            .O(N__18095),
            .I(N__18092));
    Odrv12 I__2735 (
            .O(N__18092),
            .I(M_this_map_ram_read_data_6));
    CascadeMux I__2734 (
            .O(N__18089),
            .I(N__18086));
    InMux I__2733 (
            .O(N__18086),
            .I(N__18083));
    LocalMux I__2732 (
            .O(N__18083),
            .I(N__18080));
    Odrv12 I__2731 (
            .O(N__18080),
            .I(\this_ppu.m48_i_a2_0 ));
    InMux I__2730 (
            .O(N__18077),
            .I(N__18074));
    LocalMux I__2729 (
            .O(N__18074),
            .I(N__18071));
    Span4Mux_v I__2728 (
            .O(N__18071),
            .I(N__18068));
    Span4Mux_h I__2727 (
            .O(N__18068),
            .I(N__18065));
    Sp12to4 I__2726 (
            .O(N__18065),
            .I(N__18062));
    Odrv12 I__2725 (
            .O(N__18062),
            .I(\this_spr_ram.mem_out_bus5_2 ));
    InMux I__2724 (
            .O(N__18059),
            .I(N__18056));
    LocalMux I__2723 (
            .O(N__18056),
            .I(N__18053));
    Span12Mux_v I__2722 (
            .O(N__18053),
            .I(N__18050));
    Span12Mux_v I__2721 (
            .O(N__18050),
            .I(N__18047));
    Odrv12 I__2720 (
            .O(N__18047),
            .I(\this_spr_ram.mem_out_bus1_2 ));
    InMux I__2719 (
            .O(N__18044),
            .I(N__18041));
    LocalMux I__2718 (
            .O(N__18041),
            .I(N__18038));
    Sp12to4 I__2717 (
            .O(N__18038),
            .I(N__18035));
    Span12Mux_v I__2716 (
            .O(N__18035),
            .I(N__18032));
    Odrv12 I__2715 (
            .O(N__18032),
            .I(\this_spr_ram.mem_out_bus7_2 ));
    InMux I__2714 (
            .O(N__18029),
            .I(N__18026));
    LocalMux I__2713 (
            .O(N__18026),
            .I(N__18023));
    Span4Mux_v I__2712 (
            .O(N__18023),
            .I(N__18020));
    Sp12to4 I__2711 (
            .O(N__18020),
            .I(N__18017));
    Span12Mux_h I__2710 (
            .O(N__18017),
            .I(N__18014));
    Odrv12 I__2709 (
            .O(N__18014),
            .I(\this_spr_ram.mem_out_bus3_2 ));
    InMux I__2708 (
            .O(N__18011),
            .I(N__18008));
    LocalMux I__2707 (
            .O(N__18008),
            .I(N__18005));
    Sp12to4 I__2706 (
            .O(N__18005),
            .I(N__18002));
    Span12Mux_v I__2705 (
            .O(N__18002),
            .I(N__17999));
    Span12Mux_h I__2704 (
            .O(N__17999),
            .I(N__17996));
    Odrv12 I__2703 (
            .O(N__17996),
            .I(\this_spr_ram.mem_out_bus2_2 ));
    InMux I__2702 (
            .O(N__17993),
            .I(N__17990));
    LocalMux I__2701 (
            .O(N__17990),
            .I(N__17987));
    Span12Mux_v I__2700 (
            .O(N__17987),
            .I(N__17984));
    Odrv12 I__2699 (
            .O(N__17984),
            .I(\this_spr_ram.mem_out_bus6_2 ));
    CascadeMux I__2698 (
            .O(N__17981),
            .I(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_ ));
    InMux I__2697 (
            .O(N__17978),
            .I(N__17975));
    LocalMux I__2696 (
            .O(N__17975),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ));
    InMux I__2695 (
            .O(N__17972),
            .I(N__17969));
    LocalMux I__2694 (
            .O(N__17969),
            .I(N__17966));
    Sp12to4 I__2693 (
            .O(N__17966),
            .I(N__17963));
    Span12Mux_v I__2692 (
            .O(N__17963),
            .I(N__17960));
    Span12Mux_h I__2691 (
            .O(N__17960),
            .I(N__17957));
    Odrv12 I__2690 (
            .O(N__17957),
            .I(\this_spr_ram.mem_out_bus6_1 ));
    InMux I__2689 (
            .O(N__17954),
            .I(N__17951));
    LocalMux I__2688 (
            .O(N__17951),
            .I(N__17948));
    Sp12to4 I__2687 (
            .O(N__17948),
            .I(N__17945));
    Span12Mux_v I__2686 (
            .O(N__17945),
            .I(N__17942));
    Span12Mux_h I__2685 (
            .O(N__17942),
            .I(N__17939));
    Odrv12 I__2684 (
            .O(N__17939),
            .I(\this_spr_ram.mem_out_bus2_1 ));
    InMux I__2683 (
            .O(N__17936),
            .I(N__17933));
    LocalMux I__2682 (
            .O(N__17933),
            .I(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ));
    InMux I__2681 (
            .O(N__17930),
            .I(N__17927));
    LocalMux I__2680 (
            .O(N__17927),
            .I(N__17924));
    Span4Mux_h I__2679 (
            .O(N__17924),
            .I(N__17921));
    Sp12to4 I__2678 (
            .O(N__17921),
            .I(N__17918));
    Odrv12 I__2677 (
            .O(N__17918),
            .I(\this_spr_ram.mem_out_bus4_3 ));
    InMux I__2676 (
            .O(N__17915),
            .I(N__17912));
    LocalMux I__2675 (
            .O(N__17912),
            .I(N__17909));
    Span12Mux_v I__2674 (
            .O(N__17909),
            .I(N__17906));
    Odrv12 I__2673 (
            .O(N__17906),
            .I(\this_spr_ram.mem_out_bus0_3 ));
    InMux I__2672 (
            .O(N__17903),
            .I(N__17900));
    LocalMux I__2671 (
            .O(N__17900),
            .I(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ));
    CascadeMux I__2670 (
            .O(N__17897),
            .I(N__17893));
    InMux I__2669 (
            .O(N__17896),
            .I(N__17889));
    InMux I__2668 (
            .O(N__17893),
            .I(N__17886));
    InMux I__2667 (
            .O(N__17892),
            .I(N__17881));
    LocalMux I__2666 (
            .O(N__17889),
            .I(N__17877));
    LocalMux I__2665 (
            .O(N__17886),
            .I(N__17874));
    InMux I__2664 (
            .O(N__17885),
            .I(N__17869));
    InMux I__2663 (
            .O(N__17884),
            .I(N__17869));
    LocalMux I__2662 (
            .O(N__17881),
            .I(N__17866));
    InMux I__2661 (
            .O(N__17880),
            .I(N__17863));
    Span4Mux_v I__2660 (
            .O(N__17877),
            .I(N__17860));
    Odrv4 I__2659 (
            .O(N__17874),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__2658 (
            .O(N__17869),
            .I(M_this_ppu_vram_addr_3));
    Odrv12 I__2657 (
            .O(N__17866),
            .I(M_this_ppu_vram_addr_3));
    LocalMux I__2656 (
            .O(N__17863),
            .I(M_this_ppu_vram_addr_3));
    Odrv4 I__2655 (
            .O(N__17860),
            .I(M_this_ppu_vram_addr_3));
    CascadeMux I__2654 (
            .O(N__17849),
            .I(\this_vga_signals.N_22_0_cascade_ ));
    InMux I__2653 (
            .O(N__17846),
            .I(N__17843));
    LocalMux I__2652 (
            .O(N__17843),
            .I(N__17840));
    Span4Mux_h I__2651 (
            .O(N__17840),
            .I(N__17837));
    Span4Mux_v I__2650 (
            .O(N__17837),
            .I(N__17834));
    Odrv4 I__2649 (
            .O(N__17834),
            .I(N_856_i));
    InMux I__2648 (
            .O(N__17831),
            .I(N__17828));
    LocalMux I__2647 (
            .O(N__17828),
            .I(N__17825));
    Span4Mux_v I__2646 (
            .O(N__17825),
            .I(N__17822));
    Span4Mux_h I__2645 (
            .O(N__17822),
            .I(N__17819));
    Sp12to4 I__2644 (
            .O(N__17819),
            .I(N__17816));
    Odrv12 I__2643 (
            .O(N__17816),
            .I(\this_spr_ram.mem_out_bus5_3 ));
    InMux I__2642 (
            .O(N__17813),
            .I(N__17810));
    LocalMux I__2641 (
            .O(N__17810),
            .I(N__17807));
    Span12Mux_h I__2640 (
            .O(N__17807),
            .I(N__17804));
    Span12Mux_v I__2639 (
            .O(N__17804),
            .I(N__17801));
    Odrv12 I__2638 (
            .O(N__17801),
            .I(\this_spr_ram.mem_out_bus1_3 ));
    CascadeMux I__2637 (
            .O(N__17798),
            .I(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_ ));
    InMux I__2636 (
            .O(N__17795),
            .I(N__17792));
    LocalMux I__2635 (
            .O(N__17792),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3 ));
    CascadeMux I__2634 (
            .O(N__17789),
            .I(M_this_spr_ram_read_data_3_cascade_));
    InMux I__2633 (
            .O(N__17786),
            .I(N__17783));
    LocalMux I__2632 (
            .O(N__17783),
            .I(N__17780));
    Span12Mux_s11_h I__2631 (
            .O(N__17780),
            .I(N__17777));
    Odrv12 I__2630 (
            .O(N__17777),
            .I(N_25_0_i));
    InMux I__2629 (
            .O(N__17774),
            .I(N__17771));
    LocalMux I__2628 (
            .O(N__17771),
            .I(M_this_data_tmp_qZ0Z_23));
    InMux I__2627 (
            .O(N__17768),
            .I(N__17765));
    LocalMux I__2626 (
            .O(N__17765),
            .I(N__17762));
    Span4Mux_h I__2625 (
            .O(N__17762),
            .I(N__17759));
    Odrv4 I__2624 (
            .O(N__17759),
            .I(M_this_oam_ram_write_data_19));
    InMux I__2623 (
            .O(N__17756),
            .I(N__17753));
    LocalMux I__2622 (
            .O(N__17753),
            .I(N__17750));
    Odrv4 I__2621 (
            .O(N__17750),
            .I(M_this_oam_ram_write_data_28));
    InMux I__2620 (
            .O(N__17747),
            .I(N__17744));
    LocalMux I__2619 (
            .O(N__17744),
            .I(N__17741));
    Odrv4 I__2618 (
            .O(N__17741),
            .I(M_this_oam_ram_write_data_25));
    InMux I__2617 (
            .O(N__17738),
            .I(N__17735));
    LocalMux I__2616 (
            .O(N__17735),
            .I(N__17732));
    Span4Mux_h I__2615 (
            .O(N__17732),
            .I(N__17729));
    Sp12to4 I__2614 (
            .O(N__17729),
            .I(N__17726));
    Odrv12 I__2613 (
            .O(N__17726),
            .I(\this_spr_ram.mem_out_bus4_1 ));
    InMux I__2612 (
            .O(N__17723),
            .I(N__17720));
    LocalMux I__2611 (
            .O(N__17720),
            .I(N__17717));
    Span4Mux_h I__2610 (
            .O(N__17717),
            .I(N__17714));
    Odrv4 I__2609 (
            .O(N__17714),
            .I(\this_spr_ram.mem_out_bus0_1 ));
    InMux I__2608 (
            .O(N__17711),
            .I(N__17708));
    LocalMux I__2607 (
            .O(N__17708),
            .I(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ));
    CascadeMux I__2606 (
            .O(N__17705),
            .I(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ));
    InMux I__2605 (
            .O(N__17702),
            .I(N__17699));
    LocalMux I__2604 (
            .O(N__17699),
            .I(N__17696));
    Span4Mux_v I__2603 (
            .O(N__17696),
            .I(N__17693));
    Span4Mux_h I__2602 (
            .O(N__17693),
            .I(N__17690));
    Sp12to4 I__2601 (
            .O(N__17690),
            .I(N__17687));
    Odrv12 I__2600 (
            .O(N__17687),
            .I(\this_spr_ram.mem_out_bus5_1 ));
    InMux I__2599 (
            .O(N__17684),
            .I(N__17681));
    LocalMux I__2598 (
            .O(N__17681),
            .I(N__17678));
    Span12Mux_v I__2597 (
            .O(N__17678),
            .I(N__17675));
    Odrv12 I__2596 (
            .O(N__17675),
            .I(\this_spr_ram.mem_out_bus1_1 ));
    InMux I__2595 (
            .O(N__17672),
            .I(N__17669));
    LocalMux I__2594 (
            .O(N__17669),
            .I(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ));
    InMux I__2593 (
            .O(N__17666),
            .I(N__17663));
    LocalMux I__2592 (
            .O(N__17663),
            .I(N__17660));
    Span12Mux_v I__2591 (
            .O(N__17660),
            .I(N__17657));
    Span12Mux_v I__2590 (
            .O(N__17657),
            .I(N__17654));
    Odrv12 I__2589 (
            .O(N__17654),
            .I(\this_spr_ram.mem_out_bus7_1 ));
    InMux I__2588 (
            .O(N__17651),
            .I(N__17648));
    LocalMux I__2587 (
            .O(N__17648),
            .I(N__17645));
    Span4Mux_v I__2586 (
            .O(N__17645),
            .I(N__17642));
    Sp12to4 I__2585 (
            .O(N__17642),
            .I(N__17639));
    Span12Mux_h I__2584 (
            .O(N__17639),
            .I(N__17636));
    Odrv12 I__2583 (
            .O(N__17636),
            .I(\this_spr_ram.mem_out_bus3_1 ));
    InMux I__2582 (
            .O(N__17633),
            .I(N__17630));
    LocalMux I__2581 (
            .O(N__17630),
            .I(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ));
    InMux I__2580 (
            .O(N__17627),
            .I(N__17624));
    LocalMux I__2579 (
            .O(N__17624),
            .I(N__17621));
    Span4Mux_h I__2578 (
            .O(N__17621),
            .I(N__17618));
    Odrv4 I__2577 (
            .O(N__17618),
            .I(M_this_oam_ram_write_data_1));
    InMux I__2576 (
            .O(N__17615),
            .I(N__17612));
    LocalMux I__2575 (
            .O(N__17612),
            .I(N__17609));
    Odrv4 I__2574 (
            .O(N__17609),
            .I(M_this_data_tmp_qZ0Z_20));
    InMux I__2573 (
            .O(N__17606),
            .I(N__17603));
    LocalMux I__2572 (
            .O(N__17603),
            .I(N__17600));
    Span4Mux_h I__2571 (
            .O(N__17600),
            .I(N__17597));
    Odrv4 I__2570 (
            .O(N__17597),
            .I(M_this_oam_ram_write_data_20));
    InMux I__2569 (
            .O(N__17594),
            .I(N__17591));
    LocalMux I__2568 (
            .O(N__17591),
            .I(N__17588));
    Span4Mux_h I__2567 (
            .O(N__17588),
            .I(N__17585));
    Odrv4 I__2566 (
            .O(N__17585),
            .I(M_this_oam_ram_write_data_2));
    InMux I__2565 (
            .O(N__17582),
            .I(N__17579));
    LocalMux I__2564 (
            .O(N__17579),
            .I(M_this_data_tmp_qZ0Z_9));
    InMux I__2563 (
            .O(N__17576),
            .I(N__17573));
    LocalMux I__2562 (
            .O(N__17573),
            .I(N__17570));
    Odrv4 I__2561 (
            .O(N__17570),
            .I(M_this_oam_ram_write_data_9));
    InMux I__2560 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__2559 (
            .O(N__17564),
            .I(N__17561));
    Span4Mux_h I__2558 (
            .O(N__17561),
            .I(N__17558));
    Odrv4 I__2557 (
            .O(N__17558),
            .I(M_this_oam_ram_write_data_4));
    InMux I__2556 (
            .O(N__17555),
            .I(N__17552));
    LocalMux I__2555 (
            .O(N__17552),
            .I(M_this_data_tmp_qZ0Z_11));
    InMux I__2554 (
            .O(N__17549),
            .I(N__17546));
    LocalMux I__2553 (
            .O(N__17546),
            .I(N__17543));
    Odrv12 I__2552 (
            .O(N__17543),
            .I(M_this_oam_ram_write_data_11));
    InMux I__2551 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__2550 (
            .O(N__17537),
            .I(N__17534));
    Span4Mux_s2_v I__2549 (
            .O(N__17534),
            .I(N__17531));
    Odrv4 I__2548 (
            .O(N__17531),
            .I(M_this_data_tmp_qZ0Z_17));
    InMux I__2547 (
            .O(N__17528),
            .I(N__17525));
    LocalMux I__2546 (
            .O(N__17525),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_9 ));
    InMux I__2545 (
            .O(N__17522),
            .I(N__17519));
    LocalMux I__2544 (
            .O(N__17519),
            .I(N__17516));
    Span4Mux_h I__2543 (
            .O(N__17516),
            .I(N__17513));
    Sp12to4 I__2542 (
            .O(N__17513),
            .I(N__17509));
    InMux I__2541 (
            .O(N__17512),
            .I(N__17506));
    Odrv12 I__2540 (
            .O(N__17509),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    LocalMux I__2539 (
            .O(N__17506),
            .I(\this_ppu.M_oam_cache_read_data_16 ));
    CascadeMux I__2538 (
            .O(N__17501),
            .I(N__17498));
    InMux I__2537 (
            .O(N__17498),
            .I(N__17494));
    CascadeMux I__2536 (
            .O(N__17497),
            .I(N__17491));
    LocalMux I__2535 (
            .O(N__17494),
            .I(N__17486));
    InMux I__2534 (
            .O(N__17491),
            .I(N__17483));
    CascadeMux I__2533 (
            .O(N__17490),
            .I(N__17480));
    CascadeMux I__2532 (
            .O(N__17489),
            .I(N__17476));
    Span4Mux_s0_v I__2531 (
            .O(N__17486),
            .I(N__17470));
    LocalMux I__2530 (
            .O(N__17483),
            .I(N__17470));
    InMux I__2529 (
            .O(N__17480),
            .I(N__17467));
    CascadeMux I__2528 (
            .O(N__17479),
            .I(N__17464));
    InMux I__2527 (
            .O(N__17476),
            .I(N__17459));
    CascadeMux I__2526 (
            .O(N__17475),
            .I(N__17456));
    Span4Mux_v I__2525 (
            .O(N__17470),
            .I(N__17450));
    LocalMux I__2524 (
            .O(N__17467),
            .I(N__17450));
    InMux I__2523 (
            .O(N__17464),
            .I(N__17447));
    CascadeMux I__2522 (
            .O(N__17463),
            .I(N__17444));
    CascadeMux I__2521 (
            .O(N__17462),
            .I(N__17440));
    LocalMux I__2520 (
            .O(N__17459),
            .I(N__17436));
    InMux I__2519 (
            .O(N__17456),
            .I(N__17433));
    CascadeMux I__2518 (
            .O(N__17455),
            .I(N__17430));
    Span4Mux_h I__2517 (
            .O(N__17450),
            .I(N__17423));
    LocalMux I__2516 (
            .O(N__17447),
            .I(N__17423));
    InMux I__2515 (
            .O(N__17444),
            .I(N__17420));
    CascadeMux I__2514 (
            .O(N__17443),
            .I(N__17417));
    InMux I__2513 (
            .O(N__17440),
            .I(N__17414));
    CascadeMux I__2512 (
            .O(N__17439),
            .I(N__17411));
    Span4Mux_s0_v I__2511 (
            .O(N__17436),
            .I(N__17406));
    LocalMux I__2510 (
            .O(N__17433),
            .I(N__17406));
    InMux I__2509 (
            .O(N__17430),
            .I(N__17403));
    CascadeMux I__2508 (
            .O(N__17429),
            .I(N__17400));
    CascadeMux I__2507 (
            .O(N__17428),
            .I(N__17397));
    Span4Mux_v I__2506 (
            .O(N__17423),
            .I(N__17392));
    LocalMux I__2505 (
            .O(N__17420),
            .I(N__17392));
    InMux I__2504 (
            .O(N__17417),
            .I(N__17389));
    LocalMux I__2503 (
            .O(N__17414),
            .I(N__17386));
    InMux I__2502 (
            .O(N__17411),
            .I(N__17383));
    Span4Mux_v I__2501 (
            .O(N__17406),
            .I(N__17378));
    LocalMux I__2500 (
            .O(N__17403),
            .I(N__17378));
    InMux I__2499 (
            .O(N__17400),
            .I(N__17375));
    InMux I__2498 (
            .O(N__17397),
            .I(N__17371));
    Span4Mux_v I__2497 (
            .O(N__17392),
            .I(N__17366));
    LocalMux I__2496 (
            .O(N__17389),
            .I(N__17366));
    Span4Mux_h I__2495 (
            .O(N__17386),
            .I(N__17363));
    LocalMux I__2494 (
            .O(N__17383),
            .I(N__17360));
    Span4Mux_h I__2493 (
            .O(N__17378),
            .I(N__17355));
    LocalMux I__2492 (
            .O(N__17375),
            .I(N__17355));
    CascadeMux I__2491 (
            .O(N__17374),
            .I(N__17352));
    LocalMux I__2490 (
            .O(N__17371),
            .I(N__17347));
    Span4Mux_v I__2489 (
            .O(N__17366),
            .I(N__17344));
    Span4Mux_v I__2488 (
            .O(N__17363),
            .I(N__17339));
    Span4Mux_h I__2487 (
            .O(N__17360),
            .I(N__17339));
    Span4Mux_v I__2486 (
            .O(N__17355),
            .I(N__17336));
    InMux I__2485 (
            .O(N__17352),
            .I(N__17333));
    CascadeMux I__2484 (
            .O(N__17351),
            .I(N__17330));
    CascadeMux I__2483 (
            .O(N__17350),
            .I(N__17327));
    Span12Mux_h I__2482 (
            .O(N__17347),
            .I(N__17324));
    Span4Mux_v I__2481 (
            .O(N__17344),
            .I(N__17321));
    Span4Mux_h I__2480 (
            .O(N__17339),
            .I(N__17318));
    Span4Mux_v I__2479 (
            .O(N__17336),
            .I(N__17315));
    LocalMux I__2478 (
            .O(N__17333),
            .I(N__17312));
    InMux I__2477 (
            .O(N__17330),
            .I(N__17309));
    InMux I__2476 (
            .O(N__17327),
            .I(N__17306));
    Span12Mux_v I__2475 (
            .O(N__17324),
            .I(N__17301));
    Sp12to4 I__2474 (
            .O(N__17321),
            .I(N__17301));
    Span4Mux_h I__2473 (
            .O(N__17318),
            .I(N__17298));
    Span4Mux_v I__2472 (
            .O(N__17315),
            .I(N__17295));
    Span4Mux_v I__2471 (
            .O(N__17312),
            .I(N__17288));
    LocalMux I__2470 (
            .O(N__17309),
            .I(N__17288));
    LocalMux I__2469 (
            .O(N__17306),
            .I(N__17288));
    Span12Mux_h I__2468 (
            .O(N__17301),
            .I(N__17285));
    Span4Mux_h I__2467 (
            .O(N__17298),
            .I(N__17282));
    Span4Mux_v I__2466 (
            .O(N__17295),
            .I(N__17277));
    Span4Mux_v I__2465 (
            .O(N__17288),
            .I(N__17277));
    Odrv12 I__2464 (
            .O(N__17285),
            .I(M_this_ppu_spr_addr_3));
    Odrv4 I__2463 (
            .O(N__17282),
            .I(M_this_ppu_spr_addr_3));
    Odrv4 I__2462 (
            .O(N__17277),
            .I(M_this_ppu_spr_addr_3));
    CascadeMux I__2461 (
            .O(N__17270),
            .I(N__17267));
    InMux I__2460 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__2459 (
            .O(N__17264),
            .I(N__17260));
    InMux I__2458 (
            .O(N__17263),
            .I(N__17255));
    Span4Mux_h I__2457 (
            .O(N__17260),
            .I(N__17252));
    InMux I__2456 (
            .O(N__17259),
            .I(N__17247));
    InMux I__2455 (
            .O(N__17258),
            .I(N__17247));
    LocalMux I__2454 (
            .O(N__17255),
            .I(N__17244));
    Span4Mux_v I__2453 (
            .O(N__17252),
            .I(N__17241));
    LocalMux I__2452 (
            .O(N__17247),
            .I(N__17238));
    Odrv4 I__2451 (
            .O(N__17244),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv4 I__2450 (
            .O(N__17241),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    Odrv12 I__2449 (
            .O(N__17238),
            .I(\this_ppu.M_state_qZ0Z_2 ));
    CascadeMux I__2448 (
            .O(N__17231),
            .I(N__17228));
    CascadeBuf I__2447 (
            .O(N__17228),
            .I(N__17225));
    CascadeMux I__2446 (
            .O(N__17225),
            .I(N__17222));
    InMux I__2445 (
            .O(N__17222),
            .I(N__17219));
    LocalMux I__2444 (
            .O(N__17219),
            .I(N__17216));
    Span4Mux_h I__2443 (
            .O(N__17216),
            .I(N__17211));
    InMux I__2442 (
            .O(N__17215),
            .I(N__17206));
    InMux I__2441 (
            .O(N__17214),
            .I(N__17206));
    Span4Mux_v I__2440 (
            .O(N__17211),
            .I(N__17203));
    LocalMux I__2439 (
            .O(N__17206),
            .I(M_this_oam_address_qZ0Z_6));
    Odrv4 I__2438 (
            .O(N__17203),
            .I(M_this_oam_address_qZ0Z_6));
    CascadeMux I__2437 (
            .O(N__17198),
            .I(N__17195));
    CascadeBuf I__2436 (
            .O(N__17195),
            .I(N__17192));
    CascadeMux I__2435 (
            .O(N__17192),
            .I(N__17189));
    InMux I__2434 (
            .O(N__17189),
            .I(N__17186));
    LocalMux I__2433 (
            .O(N__17186),
            .I(N__17183));
    Span4Mux_s2_v I__2432 (
            .O(N__17183),
            .I(N__17179));
    InMux I__2431 (
            .O(N__17182),
            .I(N__17176));
    Span4Mux_v I__2430 (
            .O(N__17179),
            .I(N__17173));
    LocalMux I__2429 (
            .O(N__17176),
            .I(M_this_oam_address_qZ0Z_7));
    Odrv4 I__2428 (
            .O(N__17173),
            .I(M_this_oam_address_qZ0Z_7));
    InMux I__2427 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__2426 (
            .O(N__17165),
            .I(M_this_data_tmp_qZ0Z_12));
    InMux I__2425 (
            .O(N__17162),
            .I(N__17159));
    LocalMux I__2424 (
            .O(N__17159),
            .I(N__17156));
    Odrv4 I__2423 (
            .O(N__17156),
            .I(M_this_data_tmp_qZ0Z_15));
    InMux I__2422 (
            .O(N__17153),
            .I(N__17150));
    LocalMux I__2421 (
            .O(N__17150),
            .I(N__17147));
    Odrv4 I__2420 (
            .O(N__17147),
            .I(M_this_data_tmp_qZ0Z_13));
    InMux I__2419 (
            .O(N__17144),
            .I(N__17138));
    InMux I__2418 (
            .O(N__17143),
            .I(N__17131));
    InMux I__2417 (
            .O(N__17142),
            .I(N__17131));
    InMux I__2416 (
            .O(N__17141),
            .I(N__17131));
    LocalMux I__2415 (
            .O(N__17138),
            .I(\this_ppu.N_1210_0 ));
    LocalMux I__2414 (
            .O(N__17131),
            .I(\this_ppu.N_1210_0 ));
    InMux I__2413 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__2412 (
            .O(N__17123),
            .I(\this_ppu.un1_M_screen_x_q_c3 ));
    InMux I__2411 (
            .O(N__17120),
            .I(N__17117));
    LocalMux I__2410 (
            .O(N__17117),
            .I(N__17114));
    Odrv12 I__2409 (
            .O(N__17114),
            .I(\this_ppu.oam_cache.mem_13 ));
    InMux I__2408 (
            .O(N__17111),
            .I(N__17108));
    LocalMux I__2407 (
            .O(N__17108),
            .I(N__17105));
    Odrv4 I__2406 (
            .O(N__17105),
            .I(\this_ppu.oam_cache.mem_12 ));
    InMux I__2405 (
            .O(N__17102),
            .I(N__17099));
    LocalMux I__2404 (
            .O(N__17099),
            .I(N__17096));
    Odrv4 I__2403 (
            .O(N__17096),
            .I(\this_ppu.m13_0_a2_0_0 ));
    CascadeMux I__2402 (
            .O(N__17093),
            .I(\this_ppu.N_844_cascade_ ));
    InMux I__2401 (
            .O(N__17090),
            .I(N__17084));
    InMux I__2400 (
            .O(N__17089),
            .I(N__17084));
    LocalMux I__2399 (
            .O(N__17084),
            .I(N__17080));
    InMux I__2398 (
            .O(N__17083),
            .I(N__17077));
    Odrv4 I__2397 (
            .O(N__17080),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    LocalMux I__2396 (
            .O(N__17077),
            .I(\this_ppu.M_state_qZ0Z_1 ));
    InMux I__2395 (
            .O(N__17072),
            .I(N__17068));
    InMux I__2394 (
            .O(N__17071),
            .I(N__17065));
    LocalMux I__2393 (
            .O(N__17068),
            .I(M_this_warmup_qZ0Z_1));
    LocalMux I__2392 (
            .O(N__17065),
            .I(M_this_warmup_qZ0Z_1));
    CascadeMux I__2391 (
            .O(N__17060),
            .I(N__17055));
    InMux I__2390 (
            .O(N__17059),
            .I(N__17050));
    InMux I__2389 (
            .O(N__17058),
            .I(N__17050));
    InMux I__2388 (
            .O(N__17055),
            .I(N__17047));
    LocalMux I__2387 (
            .O(N__17050),
            .I(M_this_warmup_qZ0Z_0));
    LocalMux I__2386 (
            .O(N__17047),
            .I(M_this_warmup_qZ0Z_0));
    CascadeMux I__2385 (
            .O(N__17042),
            .I(\this_ppu.N_827_0_cascade_ ));
    CascadeMux I__2384 (
            .O(N__17039),
            .I(\this_ppu.un1_M_screen_x_q_c2_cascade_ ));
    InMux I__2383 (
            .O(N__17036),
            .I(N__17033));
    LocalMux I__2382 (
            .O(N__17033),
            .I(\this_ppu.un1_M_screen_x_q_c5 ));
    CascadeMux I__2381 (
            .O(N__17030),
            .I(\this_ppu.un1_M_screen_x_q_c5_cascade_ ));
    CascadeMux I__2380 (
            .O(N__17027),
            .I(N__17024));
    InMux I__2379 (
            .O(N__17024),
            .I(N__17021));
    LocalMux I__2378 (
            .O(N__17021),
            .I(N__17018));
    Span4Mux_h I__2377 (
            .O(N__17018),
            .I(N__17013));
    InMux I__2376 (
            .O(N__17017),
            .I(N__17008));
    InMux I__2375 (
            .O(N__17016),
            .I(N__17008));
    Odrv4 I__2374 (
            .O(N__17013),
            .I(M_this_ppu_vram_addr_5));
    LocalMux I__2373 (
            .O(N__17008),
            .I(M_this_ppu_vram_addr_5));
    CascadeMux I__2372 (
            .O(N__17003),
            .I(N__17000));
    InMux I__2371 (
            .O(N__17000),
            .I(N__16997));
    LocalMux I__2370 (
            .O(N__16997),
            .I(N__16994));
    Span4Mux_h I__2369 (
            .O(N__16994),
            .I(N__16990));
    InMux I__2368 (
            .O(N__16993),
            .I(N__16987));
    Odrv4 I__2367 (
            .O(N__16990),
            .I(M_this_ppu_vram_addr_6));
    LocalMux I__2366 (
            .O(N__16987),
            .I(M_this_ppu_vram_addr_6));
    InMux I__2365 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__2364 (
            .O(N__16979),
            .I(\this_ppu.un1_M_screen_x_q_c2 ));
    CascadeMux I__2363 (
            .O(N__16976),
            .I(N__16973));
    InMux I__2362 (
            .O(N__16973),
            .I(N__16970));
    LocalMux I__2361 (
            .O(N__16970),
            .I(N__16967));
    Span4Mux_h I__2360 (
            .O(N__16967),
            .I(N__16961));
    InMux I__2359 (
            .O(N__16966),
            .I(N__16958));
    InMux I__2358 (
            .O(N__16965),
            .I(N__16953));
    InMux I__2357 (
            .O(N__16964),
            .I(N__16953));
    Odrv4 I__2356 (
            .O(N__16961),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__2355 (
            .O(N__16958),
            .I(M_this_ppu_vram_addr_1));
    LocalMux I__2354 (
            .O(N__16953),
            .I(M_this_ppu_vram_addr_1));
    CascadeMux I__2353 (
            .O(N__16946),
            .I(N__16943));
    InMux I__2352 (
            .O(N__16943),
            .I(N__16938));
    CascadeMux I__2351 (
            .O(N__16942),
            .I(N__16935));
    CascadeMux I__2350 (
            .O(N__16941),
            .I(N__16932));
    LocalMux I__2349 (
            .O(N__16938),
            .I(N__16929));
    InMux I__2348 (
            .O(N__16935),
            .I(N__16922));
    InMux I__2347 (
            .O(N__16932),
            .I(N__16922));
    Span4Mux_h I__2346 (
            .O(N__16929),
            .I(N__16919));
    InMux I__2345 (
            .O(N__16928),
            .I(N__16916));
    InMux I__2344 (
            .O(N__16927),
            .I(N__16913));
    LocalMux I__2343 (
            .O(N__16922),
            .I(M_this_ppu_vram_addr_0));
    Odrv4 I__2342 (
            .O(N__16919),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__2341 (
            .O(N__16916),
            .I(M_this_ppu_vram_addr_0));
    LocalMux I__2340 (
            .O(N__16913),
            .I(M_this_ppu_vram_addr_0));
    CascadeMux I__2339 (
            .O(N__16904),
            .I(N__16901));
    InMux I__2338 (
            .O(N__16901),
            .I(N__16897));
    CascadeMux I__2337 (
            .O(N__16900),
            .I(N__16893));
    LocalMux I__2336 (
            .O(N__16897),
            .I(N__16890));
    CascadeMux I__2335 (
            .O(N__16896),
            .I(N__16887));
    InMux I__2334 (
            .O(N__16893),
            .I(N__16884));
    Span4Mux_h I__2333 (
            .O(N__16890),
            .I(N__16880));
    InMux I__2332 (
            .O(N__16887),
            .I(N__16877));
    LocalMux I__2331 (
            .O(N__16884),
            .I(N__16874));
    InMux I__2330 (
            .O(N__16883),
            .I(N__16871));
    Odrv4 I__2329 (
            .O(N__16880),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__2328 (
            .O(N__16877),
            .I(M_this_ppu_vram_addr_2));
    Odrv4 I__2327 (
            .O(N__16874),
            .I(M_this_ppu_vram_addr_2));
    LocalMux I__2326 (
            .O(N__16871),
            .I(M_this_ppu_vram_addr_2));
    InMux I__2325 (
            .O(N__16862),
            .I(N__16855));
    InMux I__2324 (
            .O(N__16861),
            .I(N__16855));
    InMux I__2323 (
            .O(N__16860),
            .I(N__16852));
    LocalMux I__2322 (
            .O(N__16855),
            .I(\this_ppu.N_827_0 ));
    LocalMux I__2321 (
            .O(N__16852),
            .I(\this_ppu.N_827_0 ));
    CascadeMux I__2320 (
            .O(N__16847),
            .I(\this_ppu.un1_M_screen_x_q_c3_cascade_ ));
    CascadeMux I__2319 (
            .O(N__16844),
            .I(N__16841));
    InMux I__2318 (
            .O(N__16841),
            .I(N__16838));
    LocalMux I__2317 (
            .O(N__16838),
            .I(N__16835));
    Span4Mux_h I__2316 (
            .O(N__16835),
            .I(N__16830));
    InMux I__2315 (
            .O(N__16834),
            .I(N__16827));
    InMux I__2314 (
            .O(N__16833),
            .I(N__16824));
    Odrv4 I__2313 (
            .O(N__16830),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__2312 (
            .O(N__16827),
            .I(M_this_ppu_vram_addr_4));
    LocalMux I__2311 (
            .O(N__16824),
            .I(M_this_ppu_vram_addr_4));
    CascadeMux I__2310 (
            .O(N__16817),
            .I(\this_ppu.M_oam_curr_qc_0_1_cascade_ ));
    InMux I__2309 (
            .O(N__16814),
            .I(N__16811));
    LocalMux I__2308 (
            .O(N__16811),
            .I(N__16808));
    Span4Mux_h I__2307 (
            .O(N__16808),
            .I(N__16805));
    Odrv4 I__2306 (
            .O(N__16805),
            .I(\this_ppu.m35_i_a2_4 ));
    InMux I__2305 (
            .O(N__16802),
            .I(N__16799));
    LocalMux I__2304 (
            .O(N__16799),
            .I(N__16796));
    Span4Mux_s1_v I__2303 (
            .O(N__16796),
            .I(N__16793));
    Odrv4 I__2302 (
            .O(N__16793),
            .I(M_this_oam_ram_write_data_21));
    InMux I__2301 (
            .O(N__16790),
            .I(N__16787));
    LocalMux I__2300 (
            .O(N__16787),
            .I(N__16784));
    Span4Mux_s1_v I__2299 (
            .O(N__16784),
            .I(N__16781));
    Odrv4 I__2298 (
            .O(N__16781),
            .I(M_this_oam_ram_write_data_23));
    CEMux I__2297 (
            .O(N__16778),
            .I(N__16775));
    LocalMux I__2296 (
            .O(N__16775),
            .I(N__16771));
    CEMux I__2295 (
            .O(N__16774),
            .I(N__16768));
    Span4Mux_s3_v I__2294 (
            .O(N__16771),
            .I(N__16763));
    LocalMux I__2293 (
            .O(N__16768),
            .I(N__16763));
    Span4Mux_h I__2292 (
            .O(N__16763),
            .I(N__16760));
    Odrv4 I__2291 (
            .O(N__16760),
            .I(\this_spr_ram.mem_WE_12 ));
    CEMux I__2290 (
            .O(N__16757),
            .I(N__16754));
    LocalMux I__2289 (
            .O(N__16754),
            .I(N__16750));
    CEMux I__2288 (
            .O(N__16753),
            .I(N__16747));
    Span4Mux_v I__2287 (
            .O(N__16750),
            .I(N__16742));
    LocalMux I__2286 (
            .O(N__16747),
            .I(N__16742));
    Span4Mux_h I__2285 (
            .O(N__16742),
            .I(N__16739));
    Odrv4 I__2284 (
            .O(N__16739),
            .I(\this_spr_ram.mem_WE_14 ));
    InMux I__2283 (
            .O(N__16736),
            .I(N__16733));
    LocalMux I__2282 (
            .O(N__16733),
            .I(N__16730));
    Span4Mux_h I__2281 (
            .O(N__16730),
            .I(N__16727));
    Span4Mux_v I__2280 (
            .O(N__16727),
            .I(N__16724));
    Odrv4 I__2279 (
            .O(N__16724),
            .I(\this_ppu.oam_cache.mem_5 ));
    CEMux I__2278 (
            .O(N__16721),
            .I(N__16718));
    LocalMux I__2277 (
            .O(N__16718),
            .I(N__16715));
    Span4Mux_v I__2276 (
            .O(N__16715),
            .I(N__16711));
    CEMux I__2275 (
            .O(N__16714),
            .I(N__16708));
    Sp12to4 I__2274 (
            .O(N__16711),
            .I(N__16703));
    LocalMux I__2273 (
            .O(N__16708),
            .I(N__16703));
    Span12Mux_h I__2272 (
            .O(N__16703),
            .I(N__16700));
    Span12Mux_v I__2271 (
            .O(N__16700),
            .I(N__16697));
    Odrv12 I__2270 (
            .O(N__16697),
            .I(\this_spr_ram.mem_WE_0 ));
    InMux I__2269 (
            .O(N__16694),
            .I(N__16691));
    LocalMux I__2268 (
            .O(N__16691),
            .I(N__16688));
    Span4Mux_v I__2267 (
            .O(N__16688),
            .I(N__16685));
    Odrv4 I__2266 (
            .O(N__16685),
            .I(N_34_i));
    InMux I__2265 (
            .O(N__16682),
            .I(N__16679));
    LocalMux I__2264 (
            .O(N__16679),
            .I(N__16676));
    Span4Mux_v I__2263 (
            .O(N__16676),
            .I(N__16673));
    Span4Mux_h I__2262 (
            .O(N__16673),
            .I(N__16670));
    Odrv4 I__2261 (
            .O(N__16670),
            .I(\this_ppu.oam_cache.mem_14 ));
    InMux I__2260 (
            .O(N__16667),
            .I(N__16664));
    LocalMux I__2259 (
            .O(N__16664),
            .I(M_this_data_tmp_qZ0Z_8));
    InMux I__2258 (
            .O(N__16661),
            .I(N__16658));
    LocalMux I__2257 (
            .O(N__16658),
            .I(M_this_data_tmp_qZ0Z_14));
    InMux I__2256 (
            .O(N__16655),
            .I(N__16652));
    LocalMux I__2255 (
            .O(N__16652),
            .I(M_this_data_tmp_qZ0Z_10));
    InMux I__2254 (
            .O(N__16649),
            .I(N__16646));
    LocalMux I__2253 (
            .O(N__16646),
            .I(N__16643));
    Span4Mux_h I__2252 (
            .O(N__16643),
            .I(N__16640));
    Odrv4 I__2251 (
            .O(N__16640),
            .I(M_this_oam_ram_write_data_10));
    InMux I__2250 (
            .O(N__16637),
            .I(N__16634));
    LocalMux I__2249 (
            .O(N__16634),
            .I(N__16631));
    Span4Mux_v I__2248 (
            .O(N__16631),
            .I(N__16628));
    Odrv4 I__2247 (
            .O(N__16628),
            .I(M_this_oam_ram_write_data_12));
    InMux I__2246 (
            .O(N__16625),
            .I(N__16622));
    LocalMux I__2245 (
            .O(N__16622),
            .I(M_this_data_tmp_qZ0Z_7));
    InMux I__2244 (
            .O(N__16619),
            .I(N__16616));
    LocalMux I__2243 (
            .O(N__16616),
            .I(M_this_data_tmp_qZ0Z_5));
    InMux I__2242 (
            .O(N__16613),
            .I(N__16610));
    LocalMux I__2241 (
            .O(N__16610),
            .I(M_this_data_tmp_qZ0Z_22));
    InMux I__2240 (
            .O(N__16607),
            .I(N__16604));
    LocalMux I__2239 (
            .O(N__16604),
            .I(M_this_data_tmp_qZ0Z_16));
    InMux I__2238 (
            .O(N__16601),
            .I(N__16598));
    LocalMux I__2237 (
            .O(N__16598),
            .I(N__16595));
    Odrv4 I__2236 (
            .O(N__16595),
            .I(M_this_oam_ram_write_data_31));
    InMux I__2235 (
            .O(N__16592),
            .I(N__16589));
    LocalMux I__2234 (
            .O(N__16589),
            .I(M_this_warmup_qZ0Z_22));
    InMux I__2233 (
            .O(N__16586),
            .I(un1_M_this_warmup_d_cry_21));
    InMux I__2232 (
            .O(N__16583),
            .I(N__16580));
    LocalMux I__2231 (
            .O(N__16580),
            .I(M_this_warmup_qZ0Z_23));
    InMux I__2230 (
            .O(N__16577),
            .I(un1_M_this_warmup_d_cry_22));
    InMux I__2229 (
            .O(N__16574),
            .I(N__16571));
    LocalMux I__2228 (
            .O(N__16571),
            .I(M_this_warmup_qZ0Z_24));
    InMux I__2227 (
            .O(N__16568),
            .I(un1_M_this_warmup_d_cry_23));
    InMux I__2226 (
            .O(N__16565),
            .I(N__16562));
    LocalMux I__2225 (
            .O(N__16562),
            .I(M_this_warmup_qZ0Z_25));
    InMux I__2224 (
            .O(N__16559),
            .I(bfn_10_23_0_));
    InMux I__2223 (
            .O(N__16556),
            .I(N__16553));
    LocalMux I__2222 (
            .O(N__16553),
            .I(M_this_warmup_qZ0Z_26));
    InMux I__2221 (
            .O(N__16550),
            .I(un1_M_this_warmup_d_cry_25));
    InMux I__2220 (
            .O(N__16547),
            .I(N__16544));
    LocalMux I__2219 (
            .O(N__16544),
            .I(M_this_warmup_qZ0Z_27));
    InMux I__2218 (
            .O(N__16541),
            .I(un1_M_this_warmup_d_cry_26));
    InMux I__2217 (
            .O(N__16538),
            .I(un1_M_this_warmup_d_cry_27));
    InMux I__2216 (
            .O(N__16535),
            .I(N__16529));
    InMux I__2215 (
            .O(N__16534),
            .I(N__16529));
    LocalMux I__2214 (
            .O(N__16529),
            .I(M_this_warmup_qZ0Z_28));
    InMux I__2213 (
            .O(N__16526),
            .I(un1_M_this_warmup_d_cry_12));
    InMux I__2212 (
            .O(N__16523),
            .I(N__16520));
    LocalMux I__2211 (
            .O(N__16520),
            .I(M_this_warmup_qZ0Z_14));
    InMux I__2210 (
            .O(N__16517),
            .I(un1_M_this_warmup_d_cry_13));
    InMux I__2209 (
            .O(N__16514),
            .I(N__16511));
    LocalMux I__2208 (
            .O(N__16511),
            .I(M_this_warmup_qZ0Z_15));
    InMux I__2207 (
            .O(N__16508),
            .I(un1_M_this_warmup_d_cry_14));
    InMux I__2206 (
            .O(N__16505),
            .I(N__16502));
    LocalMux I__2205 (
            .O(N__16502),
            .I(M_this_warmup_qZ0Z_16));
    InMux I__2204 (
            .O(N__16499),
            .I(un1_M_this_warmup_d_cry_15));
    InMux I__2203 (
            .O(N__16496),
            .I(N__16493));
    LocalMux I__2202 (
            .O(N__16493),
            .I(M_this_warmup_qZ0Z_17));
    InMux I__2201 (
            .O(N__16490),
            .I(bfn_10_22_0_));
    InMux I__2200 (
            .O(N__16487),
            .I(N__16484));
    LocalMux I__2199 (
            .O(N__16484),
            .I(M_this_warmup_qZ0Z_18));
    InMux I__2198 (
            .O(N__16481),
            .I(un1_M_this_warmup_d_cry_17));
    InMux I__2197 (
            .O(N__16478),
            .I(N__16475));
    LocalMux I__2196 (
            .O(N__16475),
            .I(M_this_warmup_qZ0Z_19));
    InMux I__2195 (
            .O(N__16472),
            .I(un1_M_this_warmup_d_cry_18));
    InMux I__2194 (
            .O(N__16469),
            .I(N__16466));
    LocalMux I__2193 (
            .O(N__16466),
            .I(M_this_warmup_qZ0Z_20));
    InMux I__2192 (
            .O(N__16463),
            .I(un1_M_this_warmup_d_cry_19));
    InMux I__2191 (
            .O(N__16460),
            .I(N__16457));
    LocalMux I__2190 (
            .O(N__16457),
            .I(M_this_warmup_qZ0Z_21));
    InMux I__2189 (
            .O(N__16454),
            .I(un1_M_this_warmup_d_cry_20));
    InMux I__2188 (
            .O(N__16451),
            .I(N__16448));
    LocalMux I__2187 (
            .O(N__16448),
            .I(M_this_warmup_qZ0Z_5));
    InMux I__2186 (
            .O(N__16445),
            .I(un1_M_this_warmup_d_cry_4));
    InMux I__2185 (
            .O(N__16442),
            .I(N__16439));
    LocalMux I__2184 (
            .O(N__16439),
            .I(M_this_warmup_qZ0Z_6));
    InMux I__2183 (
            .O(N__16436),
            .I(un1_M_this_warmup_d_cry_5));
    InMux I__2182 (
            .O(N__16433),
            .I(N__16430));
    LocalMux I__2181 (
            .O(N__16430),
            .I(M_this_warmup_qZ0Z_7));
    InMux I__2180 (
            .O(N__16427),
            .I(un1_M_this_warmup_d_cry_6));
    InMux I__2179 (
            .O(N__16424),
            .I(N__16421));
    LocalMux I__2178 (
            .O(N__16421),
            .I(M_this_warmup_qZ0Z_8));
    InMux I__2177 (
            .O(N__16418),
            .I(un1_M_this_warmup_d_cry_7));
    InMux I__2176 (
            .O(N__16415),
            .I(N__16412));
    LocalMux I__2175 (
            .O(N__16412),
            .I(M_this_warmup_qZ0Z_9));
    InMux I__2174 (
            .O(N__16409),
            .I(bfn_10_21_0_));
    InMux I__2173 (
            .O(N__16406),
            .I(N__16403));
    LocalMux I__2172 (
            .O(N__16403),
            .I(M_this_warmup_qZ0Z_10));
    InMux I__2171 (
            .O(N__16400),
            .I(un1_M_this_warmup_d_cry_9));
    InMux I__2170 (
            .O(N__16397),
            .I(N__16394));
    LocalMux I__2169 (
            .O(N__16394),
            .I(M_this_warmup_qZ0Z_11));
    InMux I__2168 (
            .O(N__16391),
            .I(un1_M_this_warmup_d_cry_10));
    InMux I__2167 (
            .O(N__16388),
            .I(N__16385));
    LocalMux I__2166 (
            .O(N__16385),
            .I(M_this_warmup_qZ0Z_12));
    InMux I__2165 (
            .O(N__16382),
            .I(un1_M_this_warmup_d_cry_11));
    InMux I__2164 (
            .O(N__16379),
            .I(N__16376));
    LocalMux I__2163 (
            .O(N__16376),
            .I(M_this_warmup_qZ0Z_13));
    InMux I__2162 (
            .O(N__16373),
            .I(N__16370));
    LocalMux I__2161 (
            .O(N__16370),
            .I(N__16367));
    Odrv12 I__2160 (
            .O(N__16367),
            .I(\this_ppu.oam_cache.mem_10 ));
    InMux I__2159 (
            .O(N__16364),
            .I(N__16361));
    LocalMux I__2158 (
            .O(N__16361),
            .I(N__16358));
    Odrv4 I__2157 (
            .O(N__16358),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_10 ));
    CascadeMux I__2156 (
            .O(N__16355),
            .I(\this_ppu.N_836_cascade_ ));
    InMux I__2155 (
            .O(N__16352),
            .I(N__16349));
    LocalMux I__2154 (
            .O(N__16349),
            .I(N__16346));
    Span4Mux_h I__2153 (
            .O(N__16346),
            .I(N__16343));
    Odrv4 I__2152 (
            .O(N__16343),
            .I(\this_ppu.oam_cache.mem_9 ));
    InMux I__2151 (
            .O(N__16340),
            .I(N__16337));
    LocalMux I__2150 (
            .O(N__16337),
            .I(M_this_warmup_qZ0Z_2));
    InMux I__2149 (
            .O(N__16334),
            .I(un1_M_this_warmup_d_cry_1));
    InMux I__2148 (
            .O(N__16331),
            .I(N__16328));
    LocalMux I__2147 (
            .O(N__16328),
            .I(M_this_warmup_qZ0Z_3));
    InMux I__2146 (
            .O(N__16325),
            .I(un1_M_this_warmup_d_cry_2));
    InMux I__2145 (
            .O(N__16322),
            .I(N__16319));
    LocalMux I__2144 (
            .O(N__16319),
            .I(M_this_warmup_qZ0Z_4));
    InMux I__2143 (
            .O(N__16316),
            .I(un1_M_this_warmup_d_cry_3));
    InMux I__2142 (
            .O(N__16313),
            .I(N__16310));
    LocalMux I__2141 (
            .O(N__16310),
            .I(N__16307));
    Span4Mux_h I__2140 (
            .O(N__16307),
            .I(N__16303));
    InMux I__2139 (
            .O(N__16306),
            .I(N__16300));
    Odrv4 I__2138 (
            .O(N__16303),
            .I(\this_vga_signals.M_pcounter_q_i_2_0 ));
    LocalMux I__2137 (
            .O(N__16300),
            .I(\this_vga_signals.M_pcounter_q_i_2_0 ));
    InMux I__2136 (
            .O(N__16295),
            .I(N__16292));
    LocalMux I__2135 (
            .O(N__16292),
            .I(\this_vga_signals.M_pcounter_q_3_0 ));
    SRMux I__2134 (
            .O(N__16289),
            .I(N__16286));
    LocalMux I__2133 (
            .O(N__16286),
            .I(N__16282));
    SRMux I__2132 (
            .O(N__16285),
            .I(N__16279));
    Span4Mux_h I__2131 (
            .O(N__16282),
            .I(N__16275));
    LocalMux I__2130 (
            .O(N__16279),
            .I(N__16272));
    SRMux I__2129 (
            .O(N__16278),
            .I(N__16269));
    Odrv4 I__2128 (
            .O(N__16275),
            .I(\this_vga_signals.N_1188_1 ));
    Odrv4 I__2127 (
            .O(N__16272),
            .I(\this_vga_signals.N_1188_1 ));
    LocalMux I__2126 (
            .O(N__16269),
            .I(\this_vga_signals.N_1188_1 ));
    CascadeMux I__2125 (
            .O(N__16262),
            .I(\this_vga_signals.N_1188_1_cascade_ ));
    CEMux I__2124 (
            .O(N__16259),
            .I(N__16256));
    LocalMux I__2123 (
            .O(N__16256),
            .I(N__16253));
    Span4Mux_h I__2122 (
            .O(N__16253),
            .I(N__16250));
    Odrv4 I__2121 (
            .O(N__16250),
            .I(\this_vga_signals.N_933_1 ));
    InMux I__2120 (
            .O(N__16247),
            .I(N__16244));
    LocalMux I__2119 (
            .O(N__16244),
            .I(N__16238));
    InMux I__2118 (
            .O(N__16243),
            .I(N__16235));
    InMux I__2117 (
            .O(N__16242),
            .I(N__16232));
    InMux I__2116 (
            .O(N__16241),
            .I(N__16229));
    Odrv4 I__2115 (
            .O(N__16238),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__2114 (
            .O(N__16235),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__2113 (
            .O(N__16232),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    LocalMux I__2112 (
            .O(N__16229),
            .I(\this_vga_signals.M_pcounter_qZ0Z_1 ));
    CascadeMux I__2111 (
            .O(N__16220),
            .I(N__16216));
    CascadeMux I__2110 (
            .O(N__16219),
            .I(N__16212));
    InMux I__2109 (
            .O(N__16216),
            .I(N__16207));
    InMux I__2108 (
            .O(N__16215),
            .I(N__16207));
    InMux I__2107 (
            .O(N__16212),
            .I(N__16204));
    LocalMux I__2106 (
            .O(N__16207),
            .I(N__16201));
    LocalMux I__2105 (
            .O(N__16204),
            .I(N__16196));
    Span4Mux_v I__2104 (
            .O(N__16201),
            .I(N__16196));
    Odrv4 I__2103 (
            .O(N__16196),
            .I(\this_vga_signals.M_pcounter_qZ0Z_0 ));
    InMux I__2102 (
            .O(N__16193),
            .I(N__16190));
    LocalMux I__2101 (
            .O(N__16190),
            .I(N_2_0));
    InMux I__2100 (
            .O(N__16187),
            .I(N__16184));
    LocalMux I__2099 (
            .O(N__16184),
            .I(M_this_vga_signals_pixel_clk_0_0));
    CascadeMux I__2098 (
            .O(N__16181),
            .I(N_2_0_cascade_));
    InMux I__2097 (
            .O(N__16178),
            .I(N__16172));
    InMux I__2096 (
            .O(N__16177),
            .I(N__16172));
    LocalMux I__2095 (
            .O(N__16172),
            .I(N_3_0));
    InMux I__2094 (
            .O(N__16169),
            .I(N__16166));
    LocalMux I__2093 (
            .O(N__16166),
            .I(N__16161));
    InMux I__2092 (
            .O(N__16165),
            .I(N__16152));
    InMux I__2091 (
            .O(N__16164),
            .I(N__16152));
    Span4Mux_h I__2090 (
            .O(N__16161),
            .I(N__16149));
    InMux I__2089 (
            .O(N__16160),
            .I(N__16146));
    InMux I__2088 (
            .O(N__16159),
            .I(N__16139));
    InMux I__2087 (
            .O(N__16158),
            .I(N__16139));
    InMux I__2086 (
            .O(N__16157),
            .I(N__16139));
    LocalMux I__2085 (
            .O(N__16152),
            .I(N__16136));
    Odrv4 I__2084 (
            .O(N__16149),
            .I(G_462));
    LocalMux I__2083 (
            .O(N__16146),
            .I(G_462));
    LocalMux I__2082 (
            .O(N__16139),
            .I(G_462));
    Odrv4 I__2081 (
            .O(N__16136),
            .I(G_462));
    CascadeMux I__2080 (
            .O(N__16127),
            .I(N__16124));
    InMux I__2079 (
            .O(N__16124),
            .I(N__16121));
    LocalMux I__2078 (
            .O(N__16121),
            .I(\this_ppu.M_oam_cache_read_data_i_16 ));
    CascadeMux I__2077 (
            .O(N__16118),
            .I(N__16115));
    InMux I__2076 (
            .O(N__16115),
            .I(N__16112));
    LocalMux I__2075 (
            .O(N__16112),
            .I(\this_ppu.M_oam_cache_read_data_i_17 ));
    CascadeMux I__2074 (
            .O(N__16109),
            .I(N__16105));
    CascadeMux I__2073 (
            .O(N__16108),
            .I(N__16102));
    InMux I__2072 (
            .O(N__16105),
            .I(N__16098));
    InMux I__2071 (
            .O(N__16102),
            .I(N__16095));
    CascadeMux I__2070 (
            .O(N__16101),
            .I(N__16092));
    LocalMux I__2069 (
            .O(N__16098),
            .I(N__16083));
    LocalMux I__2068 (
            .O(N__16095),
            .I(N__16083));
    InMux I__2067 (
            .O(N__16092),
            .I(N__16080));
    CascadeMux I__2066 (
            .O(N__16091),
            .I(N__16077));
    CascadeMux I__2065 (
            .O(N__16090),
            .I(N__16074));
    CascadeMux I__2064 (
            .O(N__16089),
            .I(N__16069));
    CascadeMux I__2063 (
            .O(N__16088),
            .I(N__16066));
    Span4Mux_s2_v I__2062 (
            .O(N__16083),
            .I(N__16060));
    LocalMux I__2061 (
            .O(N__16080),
            .I(N__16060));
    InMux I__2060 (
            .O(N__16077),
            .I(N__16057));
    InMux I__2059 (
            .O(N__16074),
            .I(N__16054));
    CascadeMux I__2058 (
            .O(N__16073),
            .I(N__16051));
    CascadeMux I__2057 (
            .O(N__16072),
            .I(N__16048));
    InMux I__2056 (
            .O(N__16069),
            .I(N__16043));
    InMux I__2055 (
            .O(N__16066),
            .I(N__16040));
    CascadeMux I__2054 (
            .O(N__16065),
            .I(N__16037));
    Span4Mux_v I__2053 (
            .O(N__16060),
            .I(N__16032));
    LocalMux I__2052 (
            .O(N__16057),
            .I(N__16032));
    LocalMux I__2051 (
            .O(N__16054),
            .I(N__16029));
    InMux I__2050 (
            .O(N__16051),
            .I(N__16026));
    InMux I__2049 (
            .O(N__16048),
            .I(N__16023));
    CascadeMux I__2048 (
            .O(N__16047),
            .I(N__16020));
    CascadeMux I__2047 (
            .O(N__16046),
            .I(N__16017));
    LocalMux I__2046 (
            .O(N__16043),
            .I(N__16012));
    LocalMux I__2045 (
            .O(N__16040),
            .I(N__16012));
    InMux I__2044 (
            .O(N__16037),
            .I(N__16009));
    Span4Mux_v I__2043 (
            .O(N__16032),
            .I(N__15999));
    Span4Mux_h I__2042 (
            .O(N__16029),
            .I(N__15999));
    LocalMux I__2041 (
            .O(N__16026),
            .I(N__15999));
    LocalMux I__2040 (
            .O(N__16023),
            .I(N__15996));
    InMux I__2039 (
            .O(N__16020),
            .I(N__15993));
    InMux I__2038 (
            .O(N__16017),
            .I(N__15990));
    Span4Mux_s2_v I__2037 (
            .O(N__16012),
            .I(N__15985));
    LocalMux I__2036 (
            .O(N__16009),
            .I(N__15985));
    CascadeMux I__2035 (
            .O(N__16008),
            .I(N__15982));
    CascadeMux I__2034 (
            .O(N__16007),
            .I(N__15979));
    CascadeMux I__2033 (
            .O(N__16006),
            .I(N__15976));
    Span4Mux_v I__2032 (
            .O(N__15999),
            .I(N__15968));
    Span4Mux_h I__2031 (
            .O(N__15996),
            .I(N__15968));
    LocalMux I__2030 (
            .O(N__15993),
            .I(N__15968));
    LocalMux I__2029 (
            .O(N__15990),
            .I(N__15965));
    Span4Mux_v I__2028 (
            .O(N__15985),
            .I(N__15962));
    InMux I__2027 (
            .O(N__15982),
            .I(N__15959));
    InMux I__2026 (
            .O(N__15979),
            .I(N__15956));
    InMux I__2025 (
            .O(N__15976),
            .I(N__15953));
    CascadeMux I__2024 (
            .O(N__15975),
            .I(N__15950));
    Span4Mux_v I__2023 (
            .O(N__15968),
            .I(N__15947));
    Span12Mux_h I__2022 (
            .O(N__15965),
            .I(N__15940));
    Sp12to4 I__2021 (
            .O(N__15962),
            .I(N__15940));
    LocalMux I__2020 (
            .O(N__15959),
            .I(N__15940));
    LocalMux I__2019 (
            .O(N__15956),
            .I(N__15937));
    LocalMux I__2018 (
            .O(N__15953),
            .I(N__15934));
    InMux I__2017 (
            .O(N__15950),
            .I(N__15931));
    Sp12to4 I__2016 (
            .O(N__15947),
            .I(N__15928));
    Span12Mux_h I__2015 (
            .O(N__15940),
            .I(N__15925));
    Span4Mux_v I__2014 (
            .O(N__15937),
            .I(N__15918));
    Span4Mux_v I__2013 (
            .O(N__15934),
            .I(N__15918));
    LocalMux I__2012 (
            .O(N__15931),
            .I(N__15918));
    Span12Mux_h I__2011 (
            .O(N__15928),
            .I(N__15913));
    Span12Mux_v I__2010 (
            .O(N__15925),
            .I(N__15913));
    Span4Mux_v I__2009 (
            .O(N__15918),
            .I(N__15910));
    Odrv12 I__2008 (
            .O(N__15913),
            .I(M_this_ppu_spr_addr_4));
    Odrv4 I__2007 (
            .O(N__15910),
            .I(M_this_ppu_spr_addr_4));
    InMux I__2006 (
            .O(N__15905),
            .I(\this_ppu.offset_y_cry_0 ));
    InMux I__2005 (
            .O(N__15902),
            .I(N__15899));
    LocalMux I__2004 (
            .O(N__15899),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_18 ));
    InMux I__2003 (
            .O(N__15896),
            .I(\this_ppu.offset_y_cry_1 ));
    CascadeMux I__2002 (
            .O(N__15893),
            .I(N__15890));
    InMux I__2001 (
            .O(N__15890),
            .I(N__15884));
    CascadeMux I__2000 (
            .O(N__15889),
            .I(N__15881));
    CascadeMux I__1999 (
            .O(N__15888),
            .I(N__15877));
    CascadeMux I__1998 (
            .O(N__15887),
            .I(N__15874));
    LocalMux I__1997 (
            .O(N__15884),
            .I(N__15869));
    InMux I__1996 (
            .O(N__15881),
            .I(N__15866));
    CascadeMux I__1995 (
            .O(N__15880),
            .I(N__15863));
    InMux I__1994 (
            .O(N__15877),
            .I(N__15860));
    InMux I__1993 (
            .O(N__15874),
            .I(N__15857));
    CascadeMux I__1992 (
            .O(N__15873),
            .I(N__15850));
    CascadeMux I__1991 (
            .O(N__15872),
            .I(N__15847));
    Span4Mux_h I__1990 (
            .O(N__15869),
            .I(N__15841));
    LocalMux I__1989 (
            .O(N__15866),
            .I(N__15841));
    InMux I__1988 (
            .O(N__15863),
            .I(N__15838));
    LocalMux I__1987 (
            .O(N__15860),
            .I(N__15834));
    LocalMux I__1986 (
            .O(N__15857),
            .I(N__15831));
    CascadeMux I__1985 (
            .O(N__15856),
            .I(N__15828));
    CascadeMux I__1984 (
            .O(N__15855),
            .I(N__15823));
    CascadeMux I__1983 (
            .O(N__15854),
            .I(N__15819));
    CascadeMux I__1982 (
            .O(N__15853),
            .I(N__15816));
    InMux I__1981 (
            .O(N__15850),
            .I(N__15813));
    InMux I__1980 (
            .O(N__15847),
            .I(N__15810));
    CascadeMux I__1979 (
            .O(N__15846),
            .I(N__15807));
    Span4Mux_v I__1978 (
            .O(N__15841),
            .I(N__15802));
    LocalMux I__1977 (
            .O(N__15838),
            .I(N__15802));
    CascadeMux I__1976 (
            .O(N__15837),
            .I(N__15799));
    Span4Mux_h I__1975 (
            .O(N__15834),
            .I(N__15796));
    Span4Mux_v I__1974 (
            .O(N__15831),
            .I(N__15793));
    InMux I__1973 (
            .O(N__15828),
            .I(N__15790));
    CascadeMux I__1972 (
            .O(N__15827),
            .I(N__15787));
    CascadeMux I__1971 (
            .O(N__15826),
            .I(N__15784));
    InMux I__1970 (
            .O(N__15823),
            .I(N__15781));
    CascadeMux I__1969 (
            .O(N__15822),
            .I(N__15778));
    InMux I__1968 (
            .O(N__15819),
            .I(N__15775));
    InMux I__1967 (
            .O(N__15816),
            .I(N__15772));
    LocalMux I__1966 (
            .O(N__15813),
            .I(N__15769));
    LocalMux I__1965 (
            .O(N__15810),
            .I(N__15766));
    InMux I__1964 (
            .O(N__15807),
            .I(N__15763));
    Span4Mux_h I__1963 (
            .O(N__15802),
            .I(N__15760));
    InMux I__1962 (
            .O(N__15799),
            .I(N__15757));
    Span4Mux_v I__1961 (
            .O(N__15796),
            .I(N__15754));
    Span4Mux_h I__1960 (
            .O(N__15793),
            .I(N__15751));
    LocalMux I__1959 (
            .O(N__15790),
            .I(N__15748));
    InMux I__1958 (
            .O(N__15787),
            .I(N__15745));
    InMux I__1957 (
            .O(N__15784),
            .I(N__15742));
    LocalMux I__1956 (
            .O(N__15781),
            .I(N__15739));
    InMux I__1955 (
            .O(N__15778),
            .I(N__15736));
    LocalMux I__1954 (
            .O(N__15775),
            .I(N__15733));
    LocalMux I__1953 (
            .O(N__15772),
            .I(N__15730));
    Span4Mux_h I__1952 (
            .O(N__15769),
            .I(N__15727));
    Span4Mux_h I__1951 (
            .O(N__15766),
            .I(N__15724));
    LocalMux I__1950 (
            .O(N__15763),
            .I(N__15721));
    Sp12to4 I__1949 (
            .O(N__15760),
            .I(N__15718));
    LocalMux I__1948 (
            .O(N__15757),
            .I(N__15715));
    Sp12to4 I__1947 (
            .O(N__15754),
            .I(N__15708));
    Sp12to4 I__1946 (
            .O(N__15751),
            .I(N__15708));
    Span12Mux_s10_h I__1945 (
            .O(N__15748),
            .I(N__15708));
    LocalMux I__1944 (
            .O(N__15745),
            .I(N__15705));
    LocalMux I__1943 (
            .O(N__15742),
            .I(N__15702));
    Span4Mux_h I__1942 (
            .O(N__15739),
            .I(N__15699));
    LocalMux I__1941 (
            .O(N__15736),
            .I(N__15696));
    Span12Mux_h I__1940 (
            .O(N__15733),
            .I(N__15693));
    Span12Mux_s10_h I__1939 (
            .O(N__15730),
            .I(N__15690));
    Sp12to4 I__1938 (
            .O(N__15727),
            .I(N__15687));
    Span4Mux_v I__1937 (
            .O(N__15724),
            .I(N__15682));
    Span4Mux_h I__1936 (
            .O(N__15721),
            .I(N__15682));
    Span12Mux_v I__1935 (
            .O(N__15718),
            .I(N__15677));
    Span12Mux_s10_h I__1934 (
            .O(N__15715),
            .I(N__15677));
    Span12Mux_h I__1933 (
            .O(N__15708),
            .I(N__15672));
    Span12Mux_s9_h I__1932 (
            .O(N__15705),
            .I(N__15672));
    Span4Mux_h I__1931 (
            .O(N__15702),
            .I(N__15669));
    Span4Mux_v I__1930 (
            .O(N__15699),
            .I(N__15664));
    Span4Mux_h I__1929 (
            .O(N__15696),
            .I(N__15664));
    Span12Mux_v I__1928 (
            .O(N__15693),
            .I(N__15661));
    Span12Mux_h I__1927 (
            .O(N__15690),
            .I(N__15654));
    Span12Mux_s8_v I__1926 (
            .O(N__15687),
            .I(N__15654));
    Sp12to4 I__1925 (
            .O(N__15682),
            .I(N__15654));
    Span12Mux_h I__1924 (
            .O(N__15677),
            .I(N__15647));
    Span12Mux_v I__1923 (
            .O(N__15672),
            .I(N__15647));
    Sp12to4 I__1922 (
            .O(N__15669),
            .I(N__15647));
    Span4Mux_v I__1921 (
            .O(N__15664),
            .I(N__15644));
    Odrv12 I__1920 (
            .O(N__15661),
            .I(M_this_ppu_spr_addr_5));
    Odrv12 I__1919 (
            .O(N__15654),
            .I(M_this_ppu_spr_addr_5));
    Odrv12 I__1918 (
            .O(N__15647),
            .I(M_this_ppu_spr_addr_5));
    Odrv4 I__1917 (
            .O(N__15644),
            .I(M_this_ppu_spr_addr_5));
    InMux I__1916 (
            .O(N__15635),
            .I(N__15632));
    LocalMux I__1915 (
            .O(N__15632),
            .I(N__15629));
    Span4Mux_h I__1914 (
            .O(N__15629),
            .I(N__15626));
    Sp12to4 I__1913 (
            .O(N__15626),
            .I(N__15623));
    Odrv12 I__1912 (
            .O(N__15623),
            .I(\this_ppu.oam_cache.mem_4 ));
    InMux I__1911 (
            .O(N__15620),
            .I(N__15614));
    InMux I__1910 (
            .O(N__15619),
            .I(N__15614));
    LocalMux I__1909 (
            .O(N__15614),
            .I(this_pixel_clk_M_counter_q_i_1));
    InMux I__1908 (
            .O(N__15611),
            .I(N__15606));
    InMux I__1907 (
            .O(N__15610),
            .I(N__15601));
    InMux I__1906 (
            .O(N__15609),
            .I(N__15601));
    LocalMux I__1905 (
            .O(N__15606),
            .I(this_pixel_clk_M_counter_q_0));
    LocalMux I__1904 (
            .O(N__15601),
            .I(this_pixel_clk_M_counter_q_0));
    InMux I__1903 (
            .O(N__15596),
            .I(N__15593));
    LocalMux I__1902 (
            .O(N__15593),
            .I(N__15588));
    InMux I__1901 (
            .O(N__15592),
            .I(N__15585));
    CascadeMux I__1900 (
            .O(N__15591),
            .I(N__15578));
    Sp12to4 I__1899 (
            .O(N__15588),
            .I(N__15572));
    LocalMux I__1898 (
            .O(N__15585),
            .I(N__15572));
    InMux I__1897 (
            .O(N__15584),
            .I(N__15569));
    InMux I__1896 (
            .O(N__15583),
            .I(N__15560));
    InMux I__1895 (
            .O(N__15582),
            .I(N__15560));
    InMux I__1894 (
            .O(N__15581),
            .I(N__15560));
    InMux I__1893 (
            .O(N__15578),
            .I(N__15560));
    InMux I__1892 (
            .O(N__15577),
            .I(N__15556));
    Span12Mux_v I__1891 (
            .O(N__15572),
            .I(N__15549));
    LocalMux I__1890 (
            .O(N__15569),
            .I(N__15549));
    LocalMux I__1889 (
            .O(N__15560),
            .I(N__15549));
    InMux I__1888 (
            .O(N__15559),
            .I(N__15546));
    LocalMux I__1887 (
            .O(N__15556),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    Odrv12 I__1886 (
            .O(N__15549),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    LocalMux I__1885 (
            .O(N__15546),
            .I(\this_vga_signals.M_hcounter_qZ0Z_1 ));
    InMux I__1884 (
            .O(N__15539),
            .I(N__15535));
    CascadeMux I__1883 (
            .O(N__15538),
            .I(N__15532));
    LocalMux I__1882 (
            .O(N__15535),
            .I(N__15526));
    InMux I__1881 (
            .O(N__15532),
            .I(N__15523));
    InMux I__1880 (
            .O(N__15531),
            .I(N__15520));
    InMux I__1879 (
            .O(N__15530),
            .I(N__15514));
    InMux I__1878 (
            .O(N__15529),
            .I(N__15514));
    Span12Mux_v I__1877 (
            .O(N__15526),
            .I(N__15507));
    LocalMux I__1876 (
            .O(N__15523),
            .I(N__15507));
    LocalMux I__1875 (
            .O(N__15520),
            .I(N__15507));
    InMux I__1874 (
            .O(N__15519),
            .I(N__15504));
    LocalMux I__1873 (
            .O(N__15514),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    Odrv12 I__1872 (
            .O(N__15507),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    LocalMux I__1871 (
            .O(N__15504),
            .I(\this_vga_signals.M_hcounter_qZ0Z_0 ));
    CascadeMux I__1870 (
            .O(N__15497),
            .I(N_3_0_cascade_));
    InMux I__1869 (
            .O(N__15494),
            .I(N__15488));
    InMux I__1868 (
            .O(N__15493),
            .I(N__15488));
    LocalMux I__1867 (
            .O(N__15488),
            .I(N__15485));
    Odrv4 I__1866 (
            .O(N__15485),
            .I(M_this_oam_ram_read_data_20));
    InMux I__1865 (
            .O(N__15482),
            .I(N__15479));
    LocalMux I__1864 (
            .O(N__15479),
            .I(N__15476));
    Span12Mux_v I__1863 (
            .O(N__15476),
            .I(N__15473));
    Odrv12 I__1862 (
            .O(N__15473),
            .I(M_this_oam_ram_read_data_i_20));
    InMux I__1861 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__1860 (
            .O(N__15467),
            .I(M_this_oam_ram_write_data_27));
    InMux I__1859 (
            .O(N__15464),
            .I(N__15461));
    LocalMux I__1858 (
            .O(N__15461),
            .I(M_this_oam_ram_write_data_30));
    InMux I__1857 (
            .O(N__15458),
            .I(N__15455));
    LocalMux I__1856 (
            .O(N__15455),
            .I(M_this_oam_ram_write_data_17));
    InMux I__1855 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__1854 (
            .O(N__15449),
            .I(M_this_oam_ram_write_data_29));
    InMux I__1853 (
            .O(N__15446),
            .I(N__15443));
    LocalMux I__1852 (
            .O(N__15443),
            .I(M_this_oam_ram_write_data_24));
    IoInMux I__1851 (
            .O(N__15440),
            .I(N__15437));
    LocalMux I__1850 (
            .O(N__15437),
            .I(N__15432));
    IoInMux I__1849 (
            .O(N__15436),
            .I(N__15429));
    IoInMux I__1848 (
            .O(N__15435),
            .I(N__15426));
    IoSpan4Mux I__1847 (
            .O(N__15432),
            .I(N__15416));
    LocalMux I__1846 (
            .O(N__15429),
            .I(N__15416));
    LocalMux I__1845 (
            .O(N__15426),
            .I(N__15416));
    IoInMux I__1844 (
            .O(N__15425),
            .I(N__15413));
    IoInMux I__1843 (
            .O(N__15424),
            .I(N__15410));
    IoInMux I__1842 (
            .O(N__15423),
            .I(N__15405));
    IoSpan4Mux I__1841 (
            .O(N__15416),
            .I(N__15396));
    LocalMux I__1840 (
            .O(N__15413),
            .I(N__15396));
    LocalMux I__1839 (
            .O(N__15410),
            .I(N__15396));
    IoInMux I__1838 (
            .O(N__15409),
            .I(N__15393));
    IoInMux I__1837 (
            .O(N__15408),
            .I(N__15390));
    LocalMux I__1836 (
            .O(N__15405),
            .I(N__15387));
    IoInMux I__1835 (
            .O(N__15404),
            .I(N__15384));
    IoInMux I__1834 (
            .O(N__15403),
            .I(N__15381));
    IoSpan4Mux I__1833 (
            .O(N__15396),
            .I(N__15374));
    LocalMux I__1832 (
            .O(N__15393),
            .I(N__15374));
    LocalMux I__1831 (
            .O(N__15390),
            .I(N__15374));
    IoSpan4Mux I__1830 (
            .O(N__15387),
            .I(N__15365));
    LocalMux I__1829 (
            .O(N__15384),
            .I(N__15365));
    LocalMux I__1828 (
            .O(N__15381),
            .I(N__15365));
    IoSpan4Mux I__1827 (
            .O(N__15374),
            .I(N__15359));
    IoInMux I__1826 (
            .O(N__15373),
            .I(N__15356));
    IoInMux I__1825 (
            .O(N__15372),
            .I(N__15353));
    IoSpan4Mux I__1824 (
            .O(N__15365),
            .I(N__15349));
    IoInMux I__1823 (
            .O(N__15364),
            .I(N__15346));
    IoInMux I__1822 (
            .O(N__15363),
            .I(N__15343));
    IoInMux I__1821 (
            .O(N__15362),
            .I(N__15340));
    IoSpan4Mux I__1820 (
            .O(N__15359),
            .I(N__15337));
    LocalMux I__1819 (
            .O(N__15356),
            .I(N__15334));
    LocalMux I__1818 (
            .O(N__15353),
            .I(N__15331));
    IoInMux I__1817 (
            .O(N__15352),
            .I(N__15328));
    IoSpan4Mux I__1816 (
            .O(N__15349),
            .I(N__15323));
    LocalMux I__1815 (
            .O(N__15346),
            .I(N__15323));
    LocalMux I__1814 (
            .O(N__15343),
            .I(N__15320));
    LocalMux I__1813 (
            .O(N__15340),
            .I(N__15317));
    IoSpan4Mux I__1812 (
            .O(N__15337),
            .I(N__15312));
    IoSpan4Mux I__1811 (
            .O(N__15334),
            .I(N__15312));
    Span4Mux_s1_v I__1810 (
            .O(N__15331),
            .I(N__15308));
    LocalMux I__1809 (
            .O(N__15328),
            .I(N__15305));
    Span4Mux_s2_v I__1808 (
            .O(N__15323),
            .I(N__15302));
    Span4Mux_s2_v I__1807 (
            .O(N__15320),
            .I(N__15299));
    Span12Mux_s2_v I__1806 (
            .O(N__15317),
            .I(N__15296));
    Span4Mux_s2_h I__1805 (
            .O(N__15312),
            .I(N__15293));
    IoInMux I__1804 (
            .O(N__15311),
            .I(N__15290));
    Sp12to4 I__1803 (
            .O(N__15308),
            .I(N__15287));
    IoSpan4Mux I__1802 (
            .O(N__15305),
            .I(N__15284));
    Sp12to4 I__1801 (
            .O(N__15302),
            .I(N__15279));
    Sp12to4 I__1800 (
            .O(N__15299),
            .I(N__15279));
    Span12Mux_v I__1799 (
            .O(N__15296),
            .I(N__15276));
    Sp12to4 I__1798 (
            .O(N__15293),
            .I(N__15271));
    LocalMux I__1797 (
            .O(N__15290),
            .I(N__15271));
    Span12Mux_h I__1796 (
            .O(N__15287),
            .I(N__15268));
    Span4Mux_s2_h I__1795 (
            .O(N__15284),
            .I(N__15265));
    Span12Mux_h I__1794 (
            .O(N__15279),
            .I(N__15262));
    Span12Mux_v I__1793 (
            .O(N__15276),
            .I(N__15257));
    Span12Mux_s10_h I__1792 (
            .O(N__15271),
            .I(N__15257));
    Span12Mux_v I__1791 (
            .O(N__15268),
            .I(N__15252));
    Sp12to4 I__1790 (
            .O(N__15265),
            .I(N__15252));
    Span12Mux_v I__1789 (
            .O(N__15262),
            .I(N__15247));
    Span12Mux_h I__1788 (
            .O(N__15257),
            .I(N__15247));
    Span12Mux_v I__1787 (
            .O(N__15252),
            .I(N__15244));
    Odrv12 I__1786 (
            .O(N__15247),
            .I(dma_0_i));
    Odrv12 I__1785 (
            .O(N__15244),
            .I(dma_0_i));
    InMux I__1784 (
            .O(N__15239),
            .I(N__15236));
    LocalMux I__1783 (
            .O(N__15236),
            .I(N__15233));
    Span4Mux_h I__1782 (
            .O(N__15233),
            .I(N__15230));
    Sp12to4 I__1781 (
            .O(N__15230),
            .I(N__15227));
    Odrv12 I__1780 (
            .O(N__15227),
            .I(\this_ppu.oam_cache.mem_7 ));
    InMux I__1779 (
            .O(N__15224),
            .I(N__15221));
    LocalMux I__1778 (
            .O(N__15221),
            .I(N__15218));
    Span12Mux_h I__1777 (
            .O(N__15218),
            .I(N__15215));
    Odrv12 I__1776 (
            .O(N__15215),
            .I(\this_ppu.oam_cache.mem_3 ));
    InMux I__1775 (
            .O(N__15212),
            .I(N__15209));
    LocalMux I__1774 (
            .O(N__15209),
            .I(M_this_oam_ram_write_data_5));
    InMux I__1773 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__1772 (
            .O(N__15203),
            .I(N__15200));
    Odrv4 I__1771 (
            .O(N__15200),
            .I(M_this_oam_ram_write_data_7));
    InMux I__1770 (
            .O(N__15197),
            .I(N__15194));
    LocalMux I__1769 (
            .O(N__15194),
            .I(M_this_oam_ram_read_data_28));
    InMux I__1768 (
            .O(N__15191),
            .I(N__15188));
    LocalMux I__1767 (
            .O(N__15188),
            .I(N__15185));
    Span4Mux_v I__1766 (
            .O(N__15185),
            .I(N__15182));
    Span4Mux_v I__1765 (
            .O(N__15182),
            .I(N__15179));
    Odrv4 I__1764 (
            .O(N__15179),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_28 ));
    InMux I__1763 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__1762 (
            .O(N__15173),
            .I(M_this_oam_ram_read_data_29));
    InMux I__1761 (
            .O(N__15170),
            .I(N__15167));
    LocalMux I__1760 (
            .O(N__15167),
            .I(N__15164));
    Sp12to4 I__1759 (
            .O(N__15164),
            .I(N__15161));
    Odrv12 I__1758 (
            .O(N__15161),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_29 ));
    InMux I__1757 (
            .O(N__15158),
            .I(N__15155));
    LocalMux I__1756 (
            .O(N__15155),
            .I(N__15152));
    Odrv4 I__1755 (
            .O(N__15152),
            .I(M_this_oam_ram_write_data_16));
    InMux I__1754 (
            .O(N__15149),
            .I(N__15146));
    LocalMux I__1753 (
            .O(N__15146),
            .I(N__15143));
    Odrv4 I__1752 (
            .O(N__15143),
            .I(M_this_oam_ram_write_data_22));
    InMux I__1751 (
            .O(N__15140),
            .I(N__15137));
    LocalMux I__1750 (
            .O(N__15137),
            .I(N__15134));
    Span12Mux_s8_h I__1749 (
            .O(N__15134),
            .I(N__15131));
    Odrv12 I__1748 (
            .O(N__15131),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_19 ));
    InMux I__1747 (
            .O(N__15128),
            .I(N__15122));
    InMux I__1746 (
            .O(N__15127),
            .I(N__15122));
    LocalMux I__1745 (
            .O(N__15122),
            .I(N__15119));
    Odrv4 I__1744 (
            .O(N__15119),
            .I(M_this_oam_ram_read_data_19));
    InMux I__1743 (
            .O(N__15116),
            .I(N__15113));
    LocalMux I__1742 (
            .O(N__15113),
            .I(N__15110));
    Span4Mux_v I__1741 (
            .O(N__15110),
            .I(N__15107));
    Span4Mux_v I__1740 (
            .O(N__15107),
            .I(N__15104));
    Odrv4 I__1739 (
            .O(N__15104),
            .I(M_this_oam_ram_read_data_i_19));
    InMux I__1738 (
            .O(N__15101),
            .I(N__15098));
    LocalMux I__1737 (
            .O(N__15098),
            .I(N__15095));
    Span4Mux_v I__1736 (
            .O(N__15095),
            .I(N__15092));
    Span4Mux_v I__1735 (
            .O(N__15092),
            .I(N__15089));
    Odrv4 I__1734 (
            .O(N__15089),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_20 ));
    InMux I__1733 (
            .O(N__15086),
            .I(N__15083));
    LocalMux I__1732 (
            .O(N__15083),
            .I(M_this_oam_ram_write_data_13));
    InMux I__1731 (
            .O(N__15080),
            .I(N__15077));
    LocalMux I__1730 (
            .O(N__15077),
            .I(M_this_oam_ram_write_data_15));
    InMux I__1729 (
            .O(N__15074),
            .I(N__15071));
    LocalMux I__1728 (
            .O(N__15071),
            .I(N__15068));
    Span4Mux_s1_v I__1727 (
            .O(N__15068),
            .I(N__15065));
    Odrv4 I__1726 (
            .O(N__15065),
            .I(M_this_oam_ram_write_data_18));
    InMux I__1725 (
            .O(N__15062),
            .I(N__15059));
    LocalMux I__1724 (
            .O(N__15059),
            .I(N__15056));
    Odrv4 I__1723 (
            .O(N__15056),
            .I(M_this_oam_ram_read_data_31));
    InMux I__1722 (
            .O(N__15053),
            .I(N__15050));
    LocalMux I__1721 (
            .O(N__15050),
            .I(N__15047));
    Span4Mux_h I__1720 (
            .O(N__15047),
            .I(N__15044));
    Span4Mux_v I__1719 (
            .O(N__15044),
            .I(N__15041));
    Odrv4 I__1718 (
            .O(N__15041),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_31 ));
    InMux I__1717 (
            .O(N__15038),
            .I(N__15035));
    LocalMux I__1716 (
            .O(N__15035),
            .I(M_this_oam_ram_write_data_8));
    InMux I__1715 (
            .O(N__15032),
            .I(N__15029));
    LocalMux I__1714 (
            .O(N__15029),
            .I(N__15026));
    Odrv4 I__1713 (
            .O(N__15026),
            .I(M_this_data_tmp_qZ0Z_3));
    InMux I__1712 (
            .O(N__15023),
            .I(N__15020));
    LocalMux I__1711 (
            .O(N__15020),
            .I(M_this_oam_ram_write_data_3));
    InMux I__1710 (
            .O(N__15017),
            .I(N__15014));
    LocalMux I__1709 (
            .O(N__15014),
            .I(N__15010));
    InMux I__1708 (
            .O(N__15013),
            .I(N__15007));
    Span12Mux_h I__1707 (
            .O(N__15010),
            .I(N__15004));
    LocalMux I__1706 (
            .O(N__15007),
            .I(N__15001));
    Odrv12 I__1705 (
            .O(N__15004),
            .I(M_this_oam_ram_read_data_21));
    Odrv4 I__1704 (
            .O(N__15001),
            .I(M_this_oam_ram_read_data_21));
    InMux I__1703 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__1702 (
            .O(N__14993),
            .I(N__14990));
    Odrv12 I__1701 (
            .O(N__14990),
            .I(M_this_oam_ram_read_data_i_21));
    InMux I__1700 (
            .O(N__14987),
            .I(N__14984));
    LocalMux I__1699 (
            .O(N__14984),
            .I(N__14981));
    Odrv4 I__1698 (
            .O(N__14981),
            .I(M_this_data_tmp_qZ0Z_6));
    InMux I__1697 (
            .O(N__14978),
            .I(N__14975));
    LocalMux I__1696 (
            .O(N__14975),
            .I(M_this_oam_ram_write_data_6));
    InMux I__1695 (
            .O(N__14972),
            .I(N__14966));
    InMux I__1694 (
            .O(N__14971),
            .I(N__14966));
    LocalMux I__1693 (
            .O(N__14966),
            .I(N__14963));
    Span4Mux_v I__1692 (
            .O(N__14963),
            .I(N__14960));
    Span4Mux_v I__1691 (
            .O(N__14960),
            .I(N__14957));
    Odrv4 I__1690 (
            .O(N__14957),
            .I(M_this_oam_ram_read_data_22));
    InMux I__1689 (
            .O(N__14954),
            .I(N__14951));
    LocalMux I__1688 (
            .O(N__14951),
            .I(M_this_oam_ram_read_data_i_22));
    InMux I__1687 (
            .O(N__14948),
            .I(N__14944));
    InMux I__1686 (
            .O(N__14947),
            .I(N__14941));
    LocalMux I__1685 (
            .O(N__14944),
            .I(N__14936));
    LocalMux I__1684 (
            .O(N__14941),
            .I(N__14936));
    Span4Mux_v I__1683 (
            .O(N__14936),
            .I(N__14933));
    Span4Mux_v I__1682 (
            .O(N__14933),
            .I(N__14930));
    Odrv4 I__1681 (
            .O(N__14930),
            .I(M_this_oam_ram_read_data_23));
    InMux I__1680 (
            .O(N__14927),
            .I(N__14924));
    LocalMux I__1679 (
            .O(N__14924),
            .I(N__14921));
    Odrv4 I__1678 (
            .O(N__14921),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_23 ));
    InMux I__1677 (
            .O(N__14918),
            .I(N__14915));
    LocalMux I__1676 (
            .O(N__14915),
            .I(N__14912));
    Span4Mux_v I__1675 (
            .O(N__14912),
            .I(N__14909));
    Span4Mux_v I__1674 (
            .O(N__14909),
            .I(N__14906));
    Odrv4 I__1673 (
            .O(N__14906),
            .I(M_this_oam_ram_read_data_24));
    InMux I__1672 (
            .O(N__14903),
            .I(N__14900));
    LocalMux I__1671 (
            .O(N__14900),
            .I(N__14897));
    Span4Mux_h I__1670 (
            .O(N__14897),
            .I(N__14894));
    Odrv4 I__1669 (
            .O(N__14894),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_24 ));
    InMux I__1668 (
            .O(N__14891),
            .I(N__14888));
    LocalMux I__1667 (
            .O(N__14888),
            .I(N__14885));
    Span4Mux_v I__1666 (
            .O(N__14885),
            .I(N__14882));
    Span4Mux_v I__1665 (
            .O(N__14882),
            .I(N__14879));
    Odrv4 I__1664 (
            .O(N__14879),
            .I(M_this_oam_ram_read_data_25));
    InMux I__1663 (
            .O(N__14876),
            .I(N__14873));
    LocalMux I__1662 (
            .O(N__14873),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_25 ));
    InMux I__1661 (
            .O(N__14870),
            .I(N__14867));
    LocalMux I__1660 (
            .O(N__14867),
            .I(N__14864));
    Span4Mux_v I__1659 (
            .O(N__14864),
            .I(N__14861));
    Span4Mux_v I__1658 (
            .O(N__14861),
            .I(N__14858));
    Odrv4 I__1657 (
            .O(N__14858),
            .I(M_this_oam_ram_read_data_26));
    InMux I__1656 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__1655 (
            .O(N__14852),
            .I(N__14849));
    Odrv4 I__1654 (
            .O(N__14849),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_26 ));
    InMux I__1653 (
            .O(N__14846),
            .I(N__14843));
    LocalMux I__1652 (
            .O(N__14843),
            .I(M_this_oam_ram_write_data_14));
    InMux I__1651 (
            .O(N__14840),
            .I(N__14837));
    LocalMux I__1650 (
            .O(N__14837),
            .I(N__14834));
    Odrv4 I__1649 (
            .O(N__14834),
            .I(M_this_oam_ram_read_data_30));
    InMux I__1648 (
            .O(N__14831),
            .I(N__14828));
    LocalMux I__1647 (
            .O(N__14828),
            .I(N__14825));
    Span4Mux_h I__1646 (
            .O(N__14825),
            .I(N__14822));
    Span4Mux_v I__1645 (
            .O(N__14822),
            .I(N__14819));
    Odrv4 I__1644 (
            .O(N__14819),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_30 ));
    InMux I__1643 (
            .O(N__14816),
            .I(N__14813));
    LocalMux I__1642 (
            .O(N__14813),
            .I(\this_ppu.M_this_oam_ram_read_data_i_17 ));
    InMux I__1641 (
            .O(N__14810),
            .I(N__14807));
    LocalMux I__1640 (
            .O(N__14807),
            .I(\this_ppu.M_this_oam_ram_read_data_i_18 ));
    InMux I__1639 (
            .O(N__14804),
            .I(N__14801));
    LocalMux I__1638 (
            .O(N__14801),
            .I(\this_ppu.m28_e_i_o2_0 ));
    InMux I__1637 (
            .O(N__14798),
            .I(\this_ppu.un1_oam_data_1_cry_2 ));
    InMux I__1636 (
            .O(N__14795),
            .I(N__14792));
    LocalMux I__1635 (
            .O(N__14792),
            .I(\this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ));
    InMux I__1634 (
            .O(N__14789),
            .I(\this_ppu.un1_oam_data_1_cry_3 ));
    CascadeMux I__1633 (
            .O(N__14786),
            .I(N__14783));
    InMux I__1632 (
            .O(N__14783),
            .I(N__14780));
    LocalMux I__1631 (
            .O(N__14780),
            .I(\this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ));
    InMux I__1630 (
            .O(N__14777),
            .I(\this_ppu.un1_oam_data_1_cry_4 ));
    InMux I__1629 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__1628 (
            .O(N__14771),
            .I(\this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ));
    InMux I__1627 (
            .O(N__14768),
            .I(\this_ppu.un1_oam_data_1_cry_5 ));
    InMux I__1626 (
            .O(N__14765),
            .I(\this_ppu.un1_oam_data_1_cry_6 ));
    InMux I__1625 (
            .O(N__14762),
            .I(N__14759));
    LocalMux I__1624 (
            .O(N__14759),
            .I(\this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0 ));
    InMux I__1623 (
            .O(N__14756),
            .I(N__14753));
    LocalMux I__1622 (
            .O(N__14753),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_21 ));
    InMux I__1621 (
            .O(N__14750),
            .I(N__14747));
    LocalMux I__1620 (
            .O(N__14747),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_22 ));
    InMux I__1619 (
            .O(N__14744),
            .I(N__14741));
    LocalMux I__1618 (
            .O(N__14741),
            .I(N__14738));
    Odrv4 I__1617 (
            .O(N__14738),
            .I(\this_ppu.oam_cache.mem_18 ));
    CascadeMux I__1616 (
            .O(N__14735),
            .I(N__14732));
    CascadeBuf I__1615 (
            .O(N__14732),
            .I(N__14729));
    CascadeMux I__1614 (
            .O(N__14729),
            .I(N__14726));
    InMux I__1613 (
            .O(N__14726),
            .I(N__14723));
    LocalMux I__1612 (
            .O(N__14723),
            .I(\this_ppu.N_777_0 ));
    CascadeMux I__1611 (
            .O(N__14720),
            .I(N__14717));
    CascadeBuf I__1610 (
            .O(N__14717),
            .I(N__14714));
    CascadeMux I__1609 (
            .O(N__14714),
            .I(N__14711));
    InMux I__1608 (
            .O(N__14711),
            .I(N__14708));
    LocalMux I__1607 (
            .O(N__14708),
            .I(\this_ppu.N_776_0 ));
    CascadeMux I__1606 (
            .O(N__14705),
            .I(\this_ppu.N_932_0_cascade_ ));
    CascadeMux I__1605 (
            .O(N__14702),
            .I(\this_ppu.un1_M_state_q_7_i_0_0_cascade_ ));
    CascadeMux I__1604 (
            .O(N__14699),
            .I(N__14696));
    CascadeBuf I__1603 (
            .O(N__14696),
            .I(N__14693));
    CascadeMux I__1602 (
            .O(N__14693),
            .I(N__14690));
    InMux I__1601 (
            .O(N__14690),
            .I(N__14687));
    LocalMux I__1600 (
            .O(N__14687),
            .I(\this_ppu.N_775_0 ));
    InMux I__1599 (
            .O(N__14684),
            .I(N__14681));
    LocalMux I__1598 (
            .O(N__14681),
            .I(\this_ppu.N_932_0 ));
    InMux I__1597 (
            .O(N__14678),
            .I(N__14672));
    InMux I__1596 (
            .O(N__14677),
            .I(N__14672));
    LocalMux I__1595 (
            .O(N__14672),
            .I(N__14669));
    Span12Mux_v I__1594 (
            .O(N__14669),
            .I(N__14666));
    Odrv12 I__1593 (
            .O(N__14666),
            .I(\this_ppu.N_838_7 ));
    InMux I__1592 (
            .O(N__14663),
            .I(N__14660));
    LocalMux I__1591 (
            .O(N__14660),
            .I(\this_ppu.M_this_oam_ram_read_data_i_16 ));
    CascadeMux I__1590 (
            .O(N__14657),
            .I(\this_vga_ramdac.m16_cascade_ ));
    InMux I__1589 (
            .O(N__14654),
            .I(N__14651));
    LocalMux I__1588 (
            .O(N__14651),
            .I(N__14648));
    Span4Mux_h I__1587 (
            .O(N__14648),
            .I(N__14645));
    Span4Mux_h I__1586 (
            .O(N__14645),
            .I(N__14641));
    InMux I__1585 (
            .O(N__14644),
            .I(N__14638));
    Odrv4 I__1584 (
            .O(N__14641),
            .I(\this_vga_ramdac.N_3141_reto ));
    LocalMux I__1583 (
            .O(N__14638),
            .I(\this_vga_ramdac.N_3141_reto ));
    CascadeMux I__1582 (
            .O(N__14633),
            .I(\this_vga_ramdac.m19_cascade_ ));
    InMux I__1581 (
            .O(N__14630),
            .I(N__14627));
    LocalMux I__1580 (
            .O(N__14627),
            .I(N__14624));
    Span4Mux_v I__1579 (
            .O(N__14624),
            .I(N__14621));
    Span4Mux_h I__1578 (
            .O(N__14621),
            .I(N__14617));
    InMux I__1577 (
            .O(N__14620),
            .I(N__14614));
    Odrv4 I__1576 (
            .O(N__14617),
            .I(\this_vga_ramdac.N_3142_reto ));
    LocalMux I__1575 (
            .O(N__14614),
            .I(\this_vga_ramdac.N_3142_reto ));
    InMux I__1574 (
            .O(N__14609),
            .I(N__14599));
    InMux I__1573 (
            .O(N__14608),
            .I(N__14599));
    InMux I__1572 (
            .O(N__14607),
            .I(N__14590));
    InMux I__1571 (
            .O(N__14606),
            .I(N__14590));
    InMux I__1570 (
            .O(N__14605),
            .I(N__14590));
    InMux I__1569 (
            .O(N__14604),
            .I(N__14590));
    LocalMux I__1568 (
            .O(N__14599),
            .I(M_this_vram_read_data_0));
    LocalMux I__1567 (
            .O(N__14590),
            .I(M_this_vram_read_data_0));
    CascadeMux I__1566 (
            .O(N__14585),
            .I(N__14582));
    InMux I__1565 (
            .O(N__14582),
            .I(N__14575));
    InMux I__1564 (
            .O(N__14581),
            .I(N__14566));
    InMux I__1563 (
            .O(N__14580),
            .I(N__14566));
    InMux I__1562 (
            .O(N__14579),
            .I(N__14566));
    InMux I__1561 (
            .O(N__14578),
            .I(N__14566));
    LocalMux I__1560 (
            .O(N__14575),
            .I(M_this_vram_read_data_2));
    LocalMux I__1559 (
            .O(N__14566),
            .I(M_this_vram_read_data_2));
    CascadeMux I__1558 (
            .O(N__14561),
            .I(N__14553));
    InMux I__1557 (
            .O(N__14560),
            .I(N__14548));
    InMux I__1556 (
            .O(N__14559),
            .I(N__14548));
    InMux I__1555 (
            .O(N__14558),
            .I(N__14539));
    InMux I__1554 (
            .O(N__14557),
            .I(N__14539));
    InMux I__1553 (
            .O(N__14556),
            .I(N__14539));
    InMux I__1552 (
            .O(N__14553),
            .I(N__14539));
    LocalMux I__1551 (
            .O(N__14548),
            .I(M_this_vram_read_data_3));
    LocalMux I__1550 (
            .O(N__14539),
            .I(M_this_vram_read_data_3));
    CascadeMux I__1549 (
            .O(N__14534),
            .I(N__14527));
    CascadeMux I__1548 (
            .O(N__14533),
            .I(N__14524));
    CascadeMux I__1547 (
            .O(N__14532),
            .I(N__14521));
    InMux I__1546 (
            .O(N__14531),
            .I(N__14515));
    InMux I__1545 (
            .O(N__14530),
            .I(N__14515));
    InMux I__1544 (
            .O(N__14527),
            .I(N__14506));
    InMux I__1543 (
            .O(N__14524),
            .I(N__14506));
    InMux I__1542 (
            .O(N__14521),
            .I(N__14506));
    InMux I__1541 (
            .O(N__14520),
            .I(N__14506));
    LocalMux I__1540 (
            .O(N__14515),
            .I(M_this_vram_read_data_1));
    LocalMux I__1539 (
            .O(N__14506),
            .I(M_this_vram_read_data_1));
    InMux I__1538 (
            .O(N__14501),
            .I(N__14498));
    LocalMux I__1537 (
            .O(N__14498),
            .I(N__14495));
    Span4Mux_h I__1536 (
            .O(N__14495),
            .I(N__14492));
    Odrv4 I__1535 (
            .O(N__14492),
            .I(\this_vga_ramdac.m6 ));
    InMux I__1534 (
            .O(N__14489),
            .I(N__14486));
    LocalMux I__1533 (
            .O(N__14486),
            .I(N__14483));
    Span4Mux_h I__1532 (
            .O(N__14483),
            .I(N__14480));
    Odrv4 I__1531 (
            .O(N__14480),
            .I(\this_ppu.oam_cache.mem_17 ));
    InMux I__1530 (
            .O(N__14477),
            .I(N__14474));
    LocalMux I__1529 (
            .O(N__14474),
            .I(\this_ppu.oam_cache.M_oam_cache_read_data_17 ));
    InMux I__1528 (
            .O(N__14471),
            .I(N__14468));
    LocalMux I__1527 (
            .O(N__14468),
            .I(N__14465));
    Span4Mux_v I__1526 (
            .O(N__14465),
            .I(N__14462));
    Odrv4 I__1525 (
            .O(N__14462),
            .I(\this_ppu.oam_cache.mem_16 ));
    InMux I__1524 (
            .O(N__14459),
            .I(N__14456));
    LocalMux I__1523 (
            .O(N__14456),
            .I(\this_vga_ramdac.i2_mux_0 ));
    InMux I__1522 (
            .O(N__14453),
            .I(N__14450));
    LocalMux I__1521 (
            .O(N__14450),
            .I(N__14447));
    Span4Mux_v I__1520 (
            .O(N__14447),
            .I(N__14443));
    CascadeMux I__1519 (
            .O(N__14446),
            .I(N__14440));
    Span4Mux_h I__1518 (
            .O(N__14443),
            .I(N__14437));
    InMux I__1517 (
            .O(N__14440),
            .I(N__14434));
    Odrv4 I__1516 (
            .O(N__14437),
            .I(\this_vga_ramdac.N_3143_reto ));
    LocalMux I__1515 (
            .O(N__14434),
            .I(\this_vga_ramdac.N_3143_reto ));
    CascadeMux I__1514 (
            .O(N__14429),
            .I(\this_vga_ramdac.i2_mux_cascade_ ));
    InMux I__1513 (
            .O(N__14426),
            .I(N__14423));
    LocalMux I__1512 (
            .O(N__14423),
            .I(N__14419));
    InMux I__1511 (
            .O(N__14422),
            .I(N__14416));
    Span4Mux_h I__1510 (
            .O(N__14419),
            .I(N__14411));
    LocalMux I__1509 (
            .O(N__14416),
            .I(N__14411));
    Odrv4 I__1508 (
            .O(N__14411),
            .I(\this_vga_ramdac.N_3140_reto ));
    CascadeMux I__1507 (
            .O(N__14408),
            .I(\this_vga_ramdac.N_24_mux_cascade_ ));
    InMux I__1506 (
            .O(N__14405),
            .I(N__14402));
    LocalMux I__1505 (
            .O(N__14402),
            .I(N__14399));
    Span4Mux_h I__1504 (
            .O(N__14399),
            .I(N__14395));
    InMux I__1503 (
            .O(N__14398),
            .I(N__14392));
    Odrv4 I__1502 (
            .O(N__14395),
            .I(\this_vga_ramdac.N_3138_reto ));
    LocalMux I__1501 (
            .O(N__14392),
            .I(\this_vga_ramdac.N_3138_reto ));
    InMux I__1500 (
            .O(N__14387),
            .I(N__14384));
    LocalMux I__1499 (
            .O(N__14384),
            .I(N__14381));
    Span4Mux_h I__1498 (
            .O(N__14381),
            .I(N__14378));
    Odrv4 I__1497 (
            .O(N__14378),
            .I(\this_ppu.oam_cache.mem_6 ));
    CascadeMux I__1496 (
            .O(N__14375),
            .I(N__14371));
    InMux I__1495 (
            .O(N__14374),
            .I(N__14365));
    InMux I__1494 (
            .O(N__14371),
            .I(N__14365));
    InMux I__1493 (
            .O(N__14370),
            .I(N__14362));
    LocalMux I__1492 (
            .O(N__14365),
            .I(N__14355));
    LocalMux I__1491 (
            .O(N__14362),
            .I(N__14352));
    CascadeMux I__1490 (
            .O(N__14361),
            .I(N__14346));
    InMux I__1489 (
            .O(N__14360),
            .I(N__14342));
    InMux I__1488 (
            .O(N__14359),
            .I(N__14339));
    InMux I__1487 (
            .O(N__14358),
            .I(N__14336));
    Span4Mux_v I__1486 (
            .O(N__14355),
            .I(N__14331));
    Span4Mux_v I__1485 (
            .O(N__14352),
            .I(N__14331));
    InMux I__1484 (
            .O(N__14351),
            .I(N__14326));
    InMux I__1483 (
            .O(N__14350),
            .I(N__14326));
    InMux I__1482 (
            .O(N__14349),
            .I(N__14319));
    InMux I__1481 (
            .O(N__14346),
            .I(N__14319));
    InMux I__1480 (
            .O(N__14345),
            .I(N__14319));
    LocalMux I__1479 (
            .O(N__14342),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1478 (
            .O(N__14339),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1477 (
            .O(N__14336),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    Odrv4 I__1476 (
            .O(N__14331),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1475 (
            .O(N__14326),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    LocalMux I__1474 (
            .O(N__14319),
            .I(\this_vga_signals.M_hcounter_qZ0Z_5 ));
    CascadeMux I__1473 (
            .O(N__14306),
            .I(N__14303));
    InMux I__1472 (
            .O(N__14303),
            .I(N__14300));
    LocalMux I__1471 (
            .O(N__14300),
            .I(\this_vga_signals.M_hcounter_d7lt7_0 ));
    InMux I__1470 (
            .O(N__14297),
            .I(N__14287));
    InMux I__1469 (
            .O(N__14296),
            .I(N__14287));
    InMux I__1468 (
            .O(N__14295),
            .I(N__14287));
    InMux I__1467 (
            .O(N__14294),
            .I(N__14284));
    LocalMux I__1466 (
            .O(N__14287),
            .I(N__14280));
    LocalMux I__1465 (
            .O(N__14284),
            .I(N__14277));
    InMux I__1464 (
            .O(N__14283),
            .I(N__14269));
    Span4Mux_v I__1463 (
            .O(N__14280),
            .I(N__14264));
    Span4Mux_v I__1462 (
            .O(N__14277),
            .I(N__14264));
    InMux I__1461 (
            .O(N__14276),
            .I(N__14257));
    InMux I__1460 (
            .O(N__14275),
            .I(N__14257));
    InMux I__1459 (
            .O(N__14274),
            .I(N__14257));
    InMux I__1458 (
            .O(N__14273),
            .I(N__14252));
    InMux I__1457 (
            .O(N__14272),
            .I(N__14252));
    LocalMux I__1456 (
            .O(N__14269),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    Odrv4 I__1455 (
            .O(N__14264),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1454 (
            .O(N__14257),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    LocalMux I__1453 (
            .O(N__14252),
            .I(\this_vga_signals.M_hcounter_qZ0Z_6 ));
    CascadeMux I__1452 (
            .O(N__14243),
            .I(N__14237));
    InMux I__1451 (
            .O(N__14242),
            .I(N__14234));
    InMux I__1450 (
            .O(N__14241),
            .I(N__14231));
    InMux I__1449 (
            .O(N__14240),
            .I(N__14226));
    InMux I__1448 (
            .O(N__14237),
            .I(N__14226));
    LocalMux I__1447 (
            .O(N__14234),
            .I(N__14221));
    LocalMux I__1446 (
            .O(N__14231),
            .I(N__14221));
    LocalMux I__1445 (
            .O(N__14226),
            .I(N__14213));
    Span4Mux_v I__1444 (
            .O(N__14221),
            .I(N__14210));
    InMux I__1443 (
            .O(N__14220),
            .I(N__14205));
    InMux I__1442 (
            .O(N__14219),
            .I(N__14205));
    CascadeMux I__1441 (
            .O(N__14218),
            .I(N__14202));
    CascadeMux I__1440 (
            .O(N__14217),
            .I(N__14199));
    InMux I__1439 (
            .O(N__14216),
            .I(N__14196));
    Span4Mux_h I__1438 (
            .O(N__14213),
            .I(N__14189));
    Span4Mux_h I__1437 (
            .O(N__14210),
            .I(N__14189));
    LocalMux I__1436 (
            .O(N__14205),
            .I(N__14189));
    InMux I__1435 (
            .O(N__14202),
            .I(N__14186));
    InMux I__1434 (
            .O(N__14199),
            .I(N__14183));
    LocalMux I__1433 (
            .O(N__14196),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    Odrv4 I__1432 (
            .O(N__14189),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1431 (
            .O(N__14186),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    LocalMux I__1430 (
            .O(N__14183),
            .I(\this_vga_signals.M_hcounter_qZ0Z_9 ));
    InMux I__1429 (
            .O(N__14174),
            .I(N__14166));
    InMux I__1428 (
            .O(N__14173),
            .I(N__14166));
    InMux I__1427 (
            .O(N__14172),
            .I(N__14162));
    InMux I__1426 (
            .O(N__14171),
            .I(N__14159));
    LocalMux I__1425 (
            .O(N__14166),
            .I(N__14156));
    InMux I__1424 (
            .O(N__14165),
            .I(N__14153));
    LocalMux I__1423 (
            .O(N__14162),
            .I(N__14150));
    LocalMux I__1422 (
            .O(N__14159),
            .I(N__14146));
    Span4Mux_h I__1421 (
            .O(N__14156),
            .I(N__14141));
    LocalMux I__1420 (
            .O(N__14153),
            .I(N__14141));
    Span4Mux_v I__1419 (
            .O(N__14150),
            .I(N__14136));
    InMux I__1418 (
            .O(N__14149),
            .I(N__14133));
    Span4Mux_h I__1417 (
            .O(N__14146),
            .I(N__14130));
    Span4Mux_h I__1416 (
            .O(N__14141),
            .I(N__14127));
    InMux I__1415 (
            .O(N__14140),
            .I(N__14124));
    InMux I__1414 (
            .O(N__14139),
            .I(N__14121));
    Odrv4 I__1413 (
            .O(N__14136),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1412 (
            .O(N__14133),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1411 (
            .O(N__14130),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    Odrv4 I__1410 (
            .O(N__14127),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1409 (
            .O(N__14124),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    LocalMux I__1408 (
            .O(N__14121),
            .I(\this_vga_signals.M_hcounter_qZ0Z_8 ));
    CascadeMux I__1407 (
            .O(N__14108),
            .I(\this_vga_signals.N_864_cascade_ ));
    InMux I__1406 (
            .O(N__14105),
            .I(N__14094));
    InMux I__1405 (
            .O(N__14104),
            .I(N__14094));
    InMux I__1404 (
            .O(N__14103),
            .I(N__14094));
    InMux I__1403 (
            .O(N__14102),
            .I(N__14090));
    InMux I__1402 (
            .O(N__14101),
            .I(N__14087));
    LocalMux I__1401 (
            .O(N__14094),
            .I(N__14084));
    InMux I__1400 (
            .O(N__14093),
            .I(N__14081));
    LocalMux I__1399 (
            .O(N__14090),
            .I(N__14078));
    LocalMux I__1398 (
            .O(N__14087),
            .I(N__14074));
    Span4Mux_h I__1397 (
            .O(N__14084),
            .I(N__14069));
    LocalMux I__1396 (
            .O(N__14081),
            .I(N__14069));
    Span4Mux_v I__1395 (
            .O(N__14078),
            .I(N__14064));
    InMux I__1394 (
            .O(N__14077),
            .I(N__14061));
    Span4Mux_h I__1393 (
            .O(N__14074),
            .I(N__14058));
    Span4Mux_h I__1392 (
            .O(N__14069),
            .I(N__14055));
    InMux I__1391 (
            .O(N__14068),
            .I(N__14052));
    InMux I__1390 (
            .O(N__14067),
            .I(N__14049));
    Odrv4 I__1389 (
            .O(N__14064),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1388 (
            .O(N__14061),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1387 (
            .O(N__14058),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    Odrv4 I__1386 (
            .O(N__14055),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1385 (
            .O(N__14052),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    LocalMux I__1384 (
            .O(N__14049),
            .I(\this_vga_signals.M_hcounter_qZ0Z_7 ));
    InMux I__1383 (
            .O(N__14036),
            .I(N__14033));
    LocalMux I__1382 (
            .O(N__14033),
            .I(N__14029));
    InMux I__1381 (
            .O(N__14032),
            .I(N__14026));
    Span4Mux_v I__1380 (
            .O(N__14029),
            .I(N__14021));
    LocalMux I__1379 (
            .O(N__14026),
            .I(N__14021));
    Odrv4 I__1378 (
            .O(N__14021),
            .I(M_this_oam_ram_read_data_5));
    InMux I__1377 (
            .O(N__14018),
            .I(N__14015));
    LocalMux I__1376 (
            .O(N__14015),
            .I(N__14011));
    InMux I__1375 (
            .O(N__14014),
            .I(N__14008));
    Span4Mux_v I__1374 (
            .O(N__14011),
            .I(N__14003));
    LocalMux I__1373 (
            .O(N__14008),
            .I(N__14003));
    Odrv4 I__1372 (
            .O(N__14003),
            .I(M_this_oam_ram_read_data_2));
    CascadeMux I__1371 (
            .O(N__14000),
            .I(\this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_ ));
    InMux I__1370 (
            .O(N__13997),
            .I(N__13994));
    LocalMux I__1369 (
            .O(N__13994),
            .I(\this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4 ));
    CascadeMux I__1368 (
            .O(N__13991),
            .I(\this_ppu.m35_i_a2_3_cascade_ ));
    CascadeMux I__1367 (
            .O(N__13988),
            .I(\this_ppu.N_802_cascade_ ));
    CascadeMux I__1366 (
            .O(N__13985),
            .I(N__13980));
    CascadeMux I__1365 (
            .O(N__13984),
            .I(N__13977));
    CascadeMux I__1364 (
            .O(N__13983),
            .I(N__13974));
    InMux I__1363 (
            .O(N__13980),
            .I(N__13969));
    InMux I__1362 (
            .O(N__13977),
            .I(N__13961));
    InMux I__1361 (
            .O(N__13974),
            .I(N__13961));
    InMux I__1360 (
            .O(N__13973),
            .I(N__13961));
    InMux I__1359 (
            .O(N__13972),
            .I(N__13956));
    LocalMux I__1358 (
            .O(N__13969),
            .I(N__13953));
    InMux I__1357 (
            .O(N__13968),
            .I(N__13950));
    LocalMux I__1356 (
            .O(N__13961),
            .I(N__13947));
    InMux I__1355 (
            .O(N__13960),
            .I(N__13944));
    InMux I__1354 (
            .O(N__13959),
            .I(N__13941));
    LocalMux I__1353 (
            .O(N__13956),
            .I(N__13930));
    Span4Mux_h I__1352 (
            .O(N__13953),
            .I(N__13930));
    LocalMux I__1351 (
            .O(N__13950),
            .I(N__13930));
    Span4Mux_v I__1350 (
            .O(N__13947),
            .I(N__13930));
    LocalMux I__1349 (
            .O(N__13944),
            .I(N__13930));
    LocalMux I__1348 (
            .O(N__13941),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    Odrv4 I__1347 (
            .O(N__13930),
            .I(\this_vga_signals.M_hcounter_qZ0Z_3 ));
    InMux I__1346 (
            .O(N__13925),
            .I(N__13921));
    CascadeMux I__1345 (
            .O(N__13924),
            .I(N__13918));
    LocalMux I__1344 (
            .O(N__13921),
            .I(N__13912));
    InMux I__1343 (
            .O(N__13918),
            .I(N__13906));
    InMux I__1342 (
            .O(N__13917),
            .I(N__13906));
    InMux I__1341 (
            .O(N__13916),
            .I(N__13901));
    InMux I__1340 (
            .O(N__13915),
            .I(N__13901));
    Span4Mux_v I__1339 (
            .O(N__13912),
            .I(N__13896));
    InMux I__1338 (
            .O(N__13911),
            .I(N__13893));
    LocalMux I__1337 (
            .O(N__13906),
            .I(N__13888));
    LocalMux I__1336 (
            .O(N__13901),
            .I(N__13888));
    InMux I__1335 (
            .O(N__13900),
            .I(N__13885));
    InMux I__1334 (
            .O(N__13899),
            .I(N__13882));
    Span4Mux_h I__1333 (
            .O(N__13896),
            .I(N__13873));
    LocalMux I__1332 (
            .O(N__13893),
            .I(N__13873));
    Span4Mux_h I__1331 (
            .O(N__13888),
            .I(N__13873));
    LocalMux I__1330 (
            .O(N__13885),
            .I(N__13873));
    LocalMux I__1329 (
            .O(N__13882),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    Odrv4 I__1328 (
            .O(N__13873),
            .I(\this_vga_signals.M_hcounter_qZ0Z_2 ));
    InMux I__1327 (
            .O(N__13868),
            .I(N__13865));
    LocalMux I__1326 (
            .O(N__13865),
            .I(N__13862));
    Span4Mux_v I__1325 (
            .O(N__13862),
            .I(N__13859));
    Span4Mux_h I__1324 (
            .O(N__13859),
            .I(N__13856));
    Odrv4 I__1323 (
            .O(N__13856),
            .I(\this_vga_signals.un2_hsynclto3_1 ));
    CascadeMux I__1322 (
            .O(N__13853),
            .I(\this_vga_signals.un2_hsynclto3_1_cascade_ ));
    CascadeMux I__1321 (
            .O(N__13850),
            .I(N__13847));
    InMux I__1320 (
            .O(N__13847),
            .I(N__13841));
    InMux I__1319 (
            .O(N__13846),
            .I(N__13835));
    InMux I__1318 (
            .O(N__13845),
            .I(N__13835));
    CascadeMux I__1317 (
            .O(N__13844),
            .I(N__13832));
    LocalMux I__1316 (
            .O(N__13841),
            .I(N__13827));
    CascadeMux I__1315 (
            .O(N__13840),
            .I(N__13822));
    LocalMux I__1314 (
            .O(N__13835),
            .I(N__13818));
    InMux I__1313 (
            .O(N__13832),
            .I(N__13813));
    InMux I__1312 (
            .O(N__13831),
            .I(N__13813));
    InMux I__1311 (
            .O(N__13830),
            .I(N__13810));
    Span4Mux_v I__1310 (
            .O(N__13827),
            .I(N__13807));
    InMux I__1309 (
            .O(N__13826),
            .I(N__13804));
    InMux I__1308 (
            .O(N__13825),
            .I(N__13797));
    InMux I__1307 (
            .O(N__13822),
            .I(N__13797));
    InMux I__1306 (
            .O(N__13821),
            .I(N__13797));
    Span4Mux_v I__1305 (
            .O(N__13818),
            .I(N__13790));
    LocalMux I__1304 (
            .O(N__13813),
            .I(N__13790));
    LocalMux I__1303 (
            .O(N__13810),
            .I(N__13790));
    Odrv4 I__1302 (
            .O(N__13807),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1301 (
            .O(N__13804),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    LocalMux I__1300 (
            .O(N__13797),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    Odrv4 I__1299 (
            .O(N__13790),
            .I(\this_vga_signals.M_hcounter_qZ0Z_4 ));
    InMux I__1298 (
            .O(N__13781),
            .I(N__13778));
    LocalMux I__1297 (
            .O(N__13778),
            .I(N__13772));
    InMux I__1296 (
            .O(N__13777),
            .I(N__13769));
    InMux I__1295 (
            .O(N__13776),
            .I(N__13764));
    InMux I__1294 (
            .O(N__13775),
            .I(N__13761));
    Span4Mux_v I__1293 (
            .O(N__13772),
            .I(N__13755));
    LocalMux I__1292 (
            .O(N__13769),
            .I(N__13755));
    InMux I__1291 (
            .O(N__13768),
            .I(N__13752));
    CascadeMux I__1290 (
            .O(N__13767),
            .I(N__13749));
    LocalMux I__1289 (
            .O(N__13764),
            .I(N__13744));
    LocalMux I__1288 (
            .O(N__13761),
            .I(N__13744));
    InMux I__1287 (
            .O(N__13760),
            .I(N__13741));
    Span4Mux_v I__1286 (
            .O(N__13755),
            .I(N__13736));
    LocalMux I__1285 (
            .O(N__13752),
            .I(N__13736));
    InMux I__1284 (
            .O(N__13749),
            .I(N__13733));
    Span12Mux_v I__1283 (
            .O(N__13744),
            .I(N__13728));
    LocalMux I__1282 (
            .O(N__13741),
            .I(N__13728));
    Span4Mux_h I__1281 (
            .O(N__13736),
            .I(N__13725));
    LocalMux I__1280 (
            .O(N__13733),
            .I(N__13722));
    Odrv12 I__1279 (
            .O(N__13728),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto ));
    Odrv4 I__1278 (
            .O(N__13725),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto ));
    Odrv4 I__1277 (
            .O(N__13722),
            .I(\this_vga_ramdac.M_this_vga_ramdac_en_reto ));
    InMux I__1276 (
            .O(N__13715),
            .I(N__13712));
    LocalMux I__1275 (
            .O(N__13712),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ));
    CascadeMux I__1274 (
            .O(N__13709),
            .I(N__13706));
    CascadeBuf I__1273 (
            .O(N__13706),
            .I(N__13701));
    CascadeMux I__1272 (
            .O(N__13705),
            .I(N__13697));
    CascadeMux I__1271 (
            .O(N__13704),
            .I(N__13694));
    CascadeMux I__1270 (
            .O(N__13701),
            .I(N__13691));
    InMux I__1269 (
            .O(N__13700),
            .I(N__13688));
    InMux I__1268 (
            .O(N__13697),
            .I(N__13683));
    InMux I__1267 (
            .O(N__13694),
            .I(N__13683));
    InMux I__1266 (
            .O(N__13691),
            .I(N__13680));
    LocalMux I__1265 (
            .O(N__13688),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ));
    LocalMux I__1264 (
            .O(N__13683),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ));
    LocalMux I__1263 (
            .O(N__13680),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ));
    InMux I__1262 (
            .O(N__13673),
            .I(N__13670));
    LocalMux I__1261 (
            .O(N__13670),
            .I(\this_ppu.oam_cache.N_826_0 ));
    InMux I__1260 (
            .O(N__13667),
            .I(N__13664));
    LocalMux I__1259 (
            .O(N__13664),
            .I(N__13661));
    Span4Mux_h I__1258 (
            .O(N__13661),
            .I(N__13658));
    Odrv4 I__1257 (
            .O(N__13658),
            .I(\this_ppu.oam_cache.N_824_0 ));
    InMux I__1256 (
            .O(N__13655),
            .I(N__13652));
    LocalMux I__1255 (
            .O(N__13652),
            .I(N__13649));
    Span4Mux_h I__1254 (
            .O(N__13649),
            .I(N__13646));
    Odrv4 I__1253 (
            .O(N__13646),
            .I(\this_ppu.oam_cache.N_821_0 ));
    InMux I__1252 (
            .O(N__13643),
            .I(N__13640));
    LocalMux I__1251 (
            .O(N__13640),
            .I(N__13637));
    Span4Mux_h I__1250 (
            .O(N__13637),
            .I(N__13634));
    Odrv4 I__1249 (
            .O(N__13634),
            .I(\this_ppu.oam_cache.N_822_0 ));
    InMux I__1248 (
            .O(N__13631),
            .I(N__13628));
    LocalMux I__1247 (
            .O(N__13628),
            .I(N__13625));
    Span4Mux_v I__1246 (
            .O(N__13625),
            .I(N__13622));
    Odrv4 I__1245 (
            .O(N__13622),
            .I(\this_ppu.oam_cache.N_819_0 ));
    InMux I__1244 (
            .O(N__13619),
            .I(N__13616));
    LocalMux I__1243 (
            .O(N__13616),
            .I(N__13613));
    Span4Mux_h I__1242 (
            .O(N__13613),
            .I(N__13610));
    Span4Mux_v I__1241 (
            .O(N__13610),
            .I(N__13607));
    Odrv4 I__1240 (
            .O(N__13607),
            .I(\this_ppu.oam_cache.N_825_0 ));
    InMux I__1239 (
            .O(N__13604),
            .I(N__13601));
    LocalMux I__1238 (
            .O(N__13601),
            .I(N__13598));
    Span4Mux_v I__1237 (
            .O(N__13598),
            .I(N__13594));
    InMux I__1236 (
            .O(N__13597),
            .I(N__13591));
    Span4Mux_v I__1235 (
            .O(N__13594),
            .I(N__13586));
    LocalMux I__1234 (
            .O(N__13591),
            .I(N__13586));
    Odrv4 I__1233 (
            .O(N__13586),
            .I(M_this_oam_ram_read_data_0));
    InMux I__1232 (
            .O(N__13583),
            .I(N__13580));
    LocalMux I__1231 (
            .O(N__13580),
            .I(N__13576));
    InMux I__1230 (
            .O(N__13579),
            .I(N__13573));
    Span12Mux_s7_h I__1229 (
            .O(N__13576),
            .I(N__13570));
    LocalMux I__1228 (
            .O(N__13573),
            .I(N__13567));
    Odrv12 I__1227 (
            .O(N__13570),
            .I(M_this_oam_ram_read_data_6));
    Odrv4 I__1226 (
            .O(N__13567),
            .I(M_this_oam_ram_read_data_6));
    InMux I__1225 (
            .O(N__13562),
            .I(N__13558));
    CascadeMux I__1224 (
            .O(N__13561),
            .I(N__13555));
    LocalMux I__1223 (
            .O(N__13558),
            .I(N__13552));
    InMux I__1222 (
            .O(N__13555),
            .I(N__13549));
    Span4Mux_v I__1221 (
            .O(N__13552),
            .I(N__13544));
    LocalMux I__1220 (
            .O(N__13549),
            .I(N__13544));
    Odrv4 I__1219 (
            .O(N__13544),
            .I(M_this_oam_ram_read_data_1));
    InMux I__1218 (
            .O(N__13541),
            .I(N__13538));
    LocalMux I__1217 (
            .O(N__13538),
            .I(N__13535));
    Span4Mux_v I__1216 (
            .O(N__13535),
            .I(N__13531));
    InMux I__1215 (
            .O(N__13534),
            .I(N__13528));
    Span4Mux_v I__1214 (
            .O(N__13531),
            .I(N__13523));
    LocalMux I__1213 (
            .O(N__13528),
            .I(N__13523));
    Odrv4 I__1212 (
            .O(N__13523),
            .I(M_this_oam_ram_read_data_3));
    InMux I__1211 (
            .O(N__13520),
            .I(N__13517));
    LocalMux I__1210 (
            .O(N__13517),
            .I(N__13513));
    InMux I__1209 (
            .O(N__13516),
            .I(N__13510));
    Span4Mux_v I__1208 (
            .O(N__13513),
            .I(N__13505));
    LocalMux I__1207 (
            .O(N__13510),
            .I(N__13505));
    Odrv4 I__1206 (
            .O(N__13505),
            .I(M_this_oam_ram_read_data_7));
    InMux I__1205 (
            .O(N__13502),
            .I(N__13499));
    LocalMux I__1204 (
            .O(N__13499),
            .I(N__13495));
    InMux I__1203 (
            .O(N__13498),
            .I(N__13492));
    Span4Mux_v I__1202 (
            .O(N__13495),
            .I(N__13487));
    LocalMux I__1201 (
            .O(N__13492),
            .I(N__13487));
    Odrv4 I__1200 (
            .O(N__13487),
            .I(M_this_oam_ram_read_data_4));
    InMux I__1199 (
            .O(N__13484),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ));
    InMux I__1198 (
            .O(N__13481),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ));
    InMux I__1197 (
            .O(N__13478),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_3 ));
    InMux I__1196 (
            .O(N__13475),
            .I(N__13471));
    InMux I__1195 (
            .O(N__13474),
            .I(N__13468));
    LocalMux I__1194 (
            .O(N__13471),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ));
    LocalMux I__1193 (
            .O(N__13468),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ));
    CascadeMux I__1192 (
            .O(N__13463),
            .I(\this_ppu.m71_i_o2_0_cascade_ ));
    InMux I__1191 (
            .O(N__13460),
            .I(N__13457));
    LocalMux I__1190 (
            .O(N__13457),
            .I(\this_ppu.m71_i_o2_1 ));
    CascadeMux I__1189 (
            .O(N__13454),
            .I(N__13451));
    CascadeBuf I__1188 (
            .O(N__13451),
            .I(N__13446));
    CascadeMux I__1187 (
            .O(N__13450),
            .I(N__13443));
    CascadeMux I__1186 (
            .O(N__13449),
            .I(N__13439));
    CascadeMux I__1185 (
            .O(N__13446),
            .I(N__13436));
    InMux I__1184 (
            .O(N__13443),
            .I(N__13431));
    InMux I__1183 (
            .O(N__13442),
            .I(N__13431));
    InMux I__1182 (
            .O(N__13439),
            .I(N__13428));
    InMux I__1181 (
            .O(N__13436),
            .I(N__13425));
    LocalMux I__1180 (
            .O(N__13431),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_0 ));
    LocalMux I__1179 (
            .O(N__13428),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_0 ));
    LocalMux I__1178 (
            .O(N__13425),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_0 ));
    InMux I__1177 (
            .O(N__13418),
            .I(N__13415));
    LocalMux I__1176 (
            .O(N__13415),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ));
    CascadeMux I__1175 (
            .O(N__13412),
            .I(N__13409));
    CascadeBuf I__1174 (
            .O(N__13409),
            .I(N__13404));
    CascadeMux I__1173 (
            .O(N__13408),
            .I(N__13401));
    CascadeMux I__1172 (
            .O(N__13407),
            .I(N__13397));
    CascadeMux I__1171 (
            .O(N__13404),
            .I(N__13394));
    InMux I__1170 (
            .O(N__13401),
            .I(N__13391));
    InMux I__1169 (
            .O(N__13400),
            .I(N__13386));
    InMux I__1168 (
            .O(N__13397),
            .I(N__13386));
    InMux I__1167 (
            .O(N__13394),
            .I(N__13383));
    LocalMux I__1166 (
            .O(N__13391),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    LocalMux I__1165 (
            .O(N__13386),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    LocalMux I__1164 (
            .O(N__13383),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ));
    CascadeMux I__1163 (
            .O(N__13376),
            .I(N__13373));
    InMux I__1162 (
            .O(N__13373),
            .I(N__13370));
    LocalMux I__1161 (
            .O(N__13370),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ));
    CascadeMux I__1160 (
            .O(N__13367),
            .I(N__13364));
    CascadeBuf I__1159 (
            .O(N__13364),
            .I(N__13361));
    CascadeMux I__1158 (
            .O(N__13361),
            .I(N__13355));
    InMux I__1157 (
            .O(N__13360),
            .I(N__13352));
    InMux I__1156 (
            .O(N__13359),
            .I(N__13349));
    InMux I__1155 (
            .O(N__13358),
            .I(N__13346));
    InMux I__1154 (
            .O(N__13355),
            .I(N__13343));
    LocalMux I__1153 (
            .O(N__13352),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    LocalMux I__1152 (
            .O(N__13349),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    LocalMux I__1151 (
            .O(N__13346),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    LocalMux I__1150 (
            .O(N__13343),
            .I(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ));
    InMux I__1149 (
            .O(N__13334),
            .I(N__13331));
    LocalMux I__1148 (
            .O(N__13331),
            .I(N__13328));
    Span4Mux_v I__1147 (
            .O(N__13328),
            .I(N__13325));
    Span4Mux_v I__1146 (
            .O(N__13325),
            .I(N__13322));
    Odrv4 I__1145 (
            .O(N__13322),
            .I(M_this_oam_ram_read_data_14));
    InMux I__1144 (
            .O(N__13319),
            .I(N__13316));
    LocalMux I__1143 (
            .O(N__13316),
            .I(N__13313));
    Odrv4 I__1142 (
            .O(N__13313),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_14 ));
    InMux I__1141 (
            .O(N__13310),
            .I(N__13307));
    LocalMux I__1140 (
            .O(N__13307),
            .I(N__13304));
    Span4Mux_v I__1139 (
            .O(N__13304),
            .I(N__13301));
    Span4Mux_v I__1138 (
            .O(N__13301),
            .I(N__13298));
    Odrv4 I__1137 (
            .O(N__13298),
            .I(M_this_oam_ram_read_data_15));
    InMux I__1136 (
            .O(N__13295),
            .I(N__13292));
    LocalMux I__1135 (
            .O(N__13292),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_15 ));
    InMux I__1134 (
            .O(N__13289),
            .I(N__13286));
    LocalMux I__1133 (
            .O(N__13286),
            .I(\this_ppu.oam_cache.N_823_0 ));
    InMux I__1132 (
            .O(N__13283),
            .I(N__13280));
    LocalMux I__1131 (
            .O(N__13280),
            .I(\this_ppu.oam_cache.N_820_0 ));
    InMux I__1130 (
            .O(N__13277),
            .I(N__13274));
    LocalMux I__1129 (
            .O(N__13274),
            .I(N__13271));
    Span4Mux_v I__1128 (
            .O(N__13271),
            .I(N__13268));
    Span4Mux_v I__1127 (
            .O(N__13268),
            .I(N__13265));
    Span4Mux_v I__1126 (
            .O(N__13265),
            .I(N__13262));
    Odrv4 I__1125 (
            .O(N__13262),
            .I(M_this_oam_ram_read_data_8));
    InMux I__1124 (
            .O(N__13259),
            .I(N__13256));
    LocalMux I__1123 (
            .O(N__13256),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_8 ));
    InMux I__1122 (
            .O(N__13253),
            .I(N__13250));
    LocalMux I__1121 (
            .O(N__13250),
            .I(N__13247));
    Span4Mux_v I__1120 (
            .O(N__13247),
            .I(N__13244));
    Sp12to4 I__1119 (
            .O(N__13244),
            .I(N__13241));
    Odrv12 I__1118 (
            .O(N__13241),
            .I(M_this_oam_ram_read_data_9));
    InMux I__1117 (
            .O(N__13238),
            .I(N__13235));
    LocalMux I__1116 (
            .O(N__13235),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_9 ));
    InMux I__1115 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__1114 (
            .O(N__13229),
            .I(N__13226));
    Span12Mux_v I__1113 (
            .O(N__13226),
            .I(N__13223));
    Odrv12 I__1112 (
            .O(N__13223),
            .I(M_this_oam_ram_read_data_10));
    InMux I__1111 (
            .O(N__13220),
            .I(N__13217));
    LocalMux I__1110 (
            .O(N__13217),
            .I(\this_ppu.oam_cache.M_oam_cache_write_data_10 ));
    InMux I__1109 (
            .O(N__13214),
            .I(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ));
    InMux I__1108 (
            .O(N__13211),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_1 ));
    InMux I__1107 (
            .O(N__13208),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_2 ));
    InMux I__1106 (
            .O(N__13205),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_3 ));
    InMux I__1105 (
            .O(N__13202),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_4 ));
    InMux I__1104 (
            .O(N__13199),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_5 ));
    InMux I__1103 (
            .O(N__13196),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_6 ));
    InMux I__1102 (
            .O(N__13193),
            .I(\this_vga_signals.un1_M_hcounter_d_cry_7 ));
    InMux I__1101 (
            .O(N__13190),
            .I(bfn_7_18_0_));
    CascadeMux I__1100 (
            .O(N__13187),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ));
    InMux I__1099 (
            .O(N__13184),
            .I(N__13180));
    InMux I__1098 (
            .O(N__13183),
            .I(N__13177));
    LocalMux I__1097 (
            .O(N__13180),
            .I(\this_vga_signals.mult1_un68_sum_c3_2 ));
    LocalMux I__1096 (
            .O(N__13177),
            .I(\this_vga_signals.mult1_un68_sum_c3_2 ));
    CascadeMux I__1095 (
            .O(N__13172),
            .I(\this_vga_signals.mult1_un68_sum_c3_2_cascade_ ));
    CascadeMux I__1094 (
            .O(N__13169),
            .I(N__13166));
    InMux I__1093 (
            .O(N__13166),
            .I(N__13163));
    LocalMux I__1092 (
            .O(N__13163),
            .I(N__13160));
    Span4Mux_h I__1091 (
            .O(N__13160),
            .I(N__13157));
    Odrv4 I__1090 (
            .O(N__13157),
            .I(M_this_vga_signals_address_3));
    CascadeMux I__1089 (
            .O(N__13154),
            .I(N__13151));
    InMux I__1088 (
            .O(N__13151),
            .I(N__13148));
    LocalMux I__1087 (
            .O(N__13148),
            .I(N__13145));
    Span4Mux_h I__1086 (
            .O(N__13145),
            .I(N__13142));
    Odrv4 I__1085 (
            .O(N__13142),
            .I(M_this_vga_signals_address_5));
    InMux I__1084 (
            .O(N__13139),
            .I(N__13135));
    InMux I__1083 (
            .O(N__13138),
            .I(N__13132));
    LocalMux I__1082 (
            .O(N__13135),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    LocalMux I__1081 (
            .O(N__13132),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2 ));
    CascadeMux I__1080 (
            .O(N__13127),
            .I(N__13124));
    InMux I__1079 (
            .O(N__13124),
            .I(N__13121));
    LocalMux I__1078 (
            .O(N__13121),
            .I(N__13118));
    Span4Mux_h I__1077 (
            .O(N__13118),
            .I(N__13115));
    Odrv4 I__1076 (
            .O(N__13115),
            .I(M_this_vga_signals_address_4));
    InMux I__1075 (
            .O(N__13112),
            .I(N__13106));
    InMux I__1074 (
            .O(N__13111),
            .I(N__13099));
    InMux I__1073 (
            .O(N__13110),
            .I(N__13099));
    InMux I__1072 (
            .O(N__13109),
            .I(N__13099));
    LocalMux I__1071 (
            .O(N__13106),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ));
    LocalMux I__1070 (
            .O(N__13099),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ));
    CascadeMux I__1069 (
            .O(N__13094),
            .I(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ));
    InMux I__1068 (
            .O(N__13091),
            .I(N__13087));
    InMux I__1067 (
            .O(N__13090),
            .I(N__13084));
    LocalMux I__1066 (
            .O(N__13087),
            .I(\this_vga_signals.SUM_3 ));
    LocalMux I__1065 (
            .O(N__13084),
            .I(\this_vga_signals.SUM_3 ));
    InMux I__1064 (
            .O(N__13079),
            .I(N__13076));
    LocalMux I__1063 (
            .O(N__13076),
            .I(\this_vga_signals.mult1_un54_sum_c3_0 ));
    CascadeMux I__1062 (
            .O(N__13073),
            .I(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ));
    InMux I__1061 (
            .O(N__13070),
            .I(N__13067));
    LocalMux I__1060 (
            .O(N__13067),
            .I(\this_vga_signals.if_m1_1 ));
    InMux I__1059 (
            .O(N__13064),
            .I(N__13061));
    LocalMux I__1058 (
            .O(N__13061),
            .I(N__13057));
    CascadeMux I__1057 (
            .O(N__13060),
            .I(N__13054));
    Span4Mux_h I__1056 (
            .O(N__13057),
            .I(N__13051));
    InMux I__1055 (
            .O(N__13054),
            .I(N__13048));
    Odrv4 I__1054 (
            .O(N__13051),
            .I(\this_vga_ramdac.N_3139_reto ));
    LocalMux I__1053 (
            .O(N__13048),
            .I(\this_vga_ramdac.N_3139_reto ));
    CascadeMux I__1052 (
            .O(N__13043),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ));
    InMux I__1051 (
            .O(N__13040),
            .I(N__13030));
    InMux I__1050 (
            .O(N__13039),
            .I(N__13030));
    InMux I__1049 (
            .O(N__13038),
            .I(N__13030));
    InMux I__1048 (
            .O(N__13037),
            .I(N__13027));
    LocalMux I__1047 (
            .O(N__13030),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    LocalMux I__1046 (
            .O(N__13027),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3 ));
    CascadeMux I__1045 (
            .O(N__13022),
            .I(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ));
    CascadeMux I__1044 (
            .O(N__13019),
            .I(N__13016));
    InMux I__1043 (
            .O(N__13016),
            .I(N__13013));
    LocalMux I__1042 (
            .O(N__13013),
            .I(N__13010));
    Odrv4 I__1041 (
            .O(N__13010),
            .I(M_this_vga_signals_address_2));
    CascadeMux I__1040 (
            .O(N__13007),
            .I(\this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_ ));
    InMux I__1039 (
            .O(N__13004),
            .I(N__13001));
    LocalMux I__1038 (
            .O(N__13001),
            .I(\this_vga_signals.if_m7_0_o4_1_ns_1 ));
    CascadeMux I__1037 (
            .O(N__12998),
            .I(\this_vga_signals.SUM_3_cascade_ ));
    InMux I__1036 (
            .O(N__12995),
            .I(N__12992));
    LocalMux I__1035 (
            .O(N__12992),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_1 ));
    InMux I__1034 (
            .O(N__12989),
            .I(N__12986));
    LocalMux I__1033 (
            .O(N__12986),
            .I(\this_vga_signals.mult1_un89_sum_c3_0 ));
    CascadeMux I__1032 (
            .O(N__12983),
            .I(N__12980));
    InMux I__1031 (
            .O(N__12980),
            .I(N__12977));
    LocalMux I__1030 (
            .O(N__12977),
            .I(N__12974));
    Odrv4 I__1029 (
            .O(N__12974),
            .I(M_this_vga_signals_address_0));
    InMux I__1028 (
            .O(N__12971),
            .I(N__12967));
    InMux I__1027 (
            .O(N__12970),
            .I(N__12964));
    LocalMux I__1026 (
            .O(N__12967),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    LocalMux I__1025 (
            .O(N__12964),
            .I(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ));
    InMux I__1024 (
            .O(N__12959),
            .I(N__12956));
    LocalMux I__1023 (
            .O(N__12956),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1_2 ));
    InMux I__1022 (
            .O(N__12953),
            .I(N__12950));
    LocalMux I__1021 (
            .O(N__12950),
            .I(\this_vga_signals.un2_hsynclto6_0 ));
    CascadeMux I__1020 (
            .O(N__12947),
            .I(\this_vga_signals.un4_hsynclt7_cascade_ ));
    InMux I__1019 (
            .O(N__12944),
            .I(N__12941));
    LocalMux I__1018 (
            .O(N__12941),
            .I(\this_vga_signals.hsync_1_1 ));
    CascadeMux I__1017 (
            .O(N__12938),
            .I(\this_vga_signals.un4_hsynclt8_0_cascade_ ));
    IoInMux I__1016 (
            .O(N__12935),
            .I(N__12932));
    LocalMux I__1015 (
            .O(N__12932),
            .I(N__12929));
    Span12Mux_s2_v I__1014 (
            .O(N__12929),
            .I(N__12926));
    Span12Mux_v I__1013 (
            .O(N__12926),
            .I(N__12923));
    Odrv12 I__1012 (
            .O(N__12923),
            .I(this_vga_signals_hsync_1_i));
    IoInMux I__1011 (
            .O(N__12920),
            .I(N__12917));
    LocalMux I__1010 (
            .O(N__12917),
            .I(N__12914));
    Span4Mux_s0_v I__1009 (
            .O(N__12914),
            .I(N__12911));
    Span4Mux_v I__1008 (
            .O(N__12911),
            .I(N__12908));
    Span4Mux_v I__1007 (
            .O(N__12908),
            .I(N__12905));
    Span4Mux_v I__1006 (
            .O(N__12905),
            .I(N__12902));
    Odrv4 I__1005 (
            .O(N__12902),
            .I(this_vga_signals_hvisibility_i));
    IoInMux I__1004 (
            .O(N__12899),
            .I(N__12896));
    LocalMux I__1003 (
            .O(N__12896),
            .I(N__12893));
    Odrv12 I__1002 (
            .O(N__12893),
            .I(this_vga_signals_vvisibility_i));
    IoInMux I__1001 (
            .O(N__12890),
            .I(N__12887));
    LocalMux I__1000 (
            .O(N__12887),
            .I(N__12884));
    Span4Mux_s1_h I__999 (
            .O(N__12884),
            .I(N__12881));
    Sp12to4 I__998 (
            .O(N__12881),
            .I(N__12878));
    Span12Mux_v I__997 (
            .O(N__12878),
            .I(N__12875));
    Odrv12 I__996 (
            .O(N__12875),
            .I(rgb_c_0));
    CascadeMux I__995 (
            .O(N__12872),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_ ));
    CascadeMux I__994 (
            .O(N__12869),
            .I(\this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ));
    InMux I__993 (
            .O(N__12866),
            .I(N__12863));
    LocalMux I__992 (
            .O(N__12863),
            .I(\this_vga_signals.mult1_un89_sum_c3_1 ));
    InMux I__991 (
            .O(N__12860),
            .I(N__12854));
    InMux I__990 (
            .O(N__12859),
            .I(N__12854));
    LocalMux I__989 (
            .O(N__12854),
            .I(\this_vga_signals.mult1_un82_sum_c3_0 ));
    InMux I__988 (
            .O(N__12851),
            .I(N__12845));
    InMux I__987 (
            .O(N__12850),
            .I(N__12845));
    LocalMux I__986 (
            .O(N__12845),
            .I(\this_vga_signals.mult1_un82_sum_axbxc3_1 ));
    CascadeMux I__985 (
            .O(N__12842),
            .I(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ));
    CascadeMux I__984 (
            .O(N__12839),
            .I(N__12836));
    InMux I__983 (
            .O(N__12836),
            .I(N__12833));
    LocalMux I__982 (
            .O(N__12833),
            .I(N__12830));
    Odrv12 I__981 (
            .O(N__12830),
            .I(M_this_vga_signals_address_1));
    InMux I__980 (
            .O(N__12827),
            .I(N__12824));
    LocalMux I__979 (
            .O(N__12824),
            .I(\this_vga_signals.SUM_3_1 ));
    CascadeMux I__978 (
            .O(N__12821),
            .I(N__12818));
    InMux I__977 (
            .O(N__12818),
            .I(N__12812));
    InMux I__976 (
            .O(N__12817),
            .I(N__12812));
    LocalMux I__975 (
            .O(N__12812),
            .I(\this_vga_signals.mult1_un75_sum_axb1 ));
    IoInMux I__974 (
            .O(N__12809),
            .I(N__12806));
    LocalMux I__973 (
            .O(N__12806),
            .I(N__12803));
    IoSpan4Mux I__972 (
            .O(N__12803),
            .I(N__12800));
    IoSpan4Mux I__971 (
            .O(N__12800),
            .I(N__12797));
    Span4Mux_s1_h I__970 (
            .O(N__12797),
            .I(N__12794));
    Odrv4 I__969 (
            .O(N__12794),
            .I(rgb_c_3));
    IoInMux I__968 (
            .O(N__12791),
            .I(N__12788));
    LocalMux I__967 (
            .O(N__12788),
            .I(N__12785));
    Odrv12 I__966 (
            .O(N__12785),
            .I(rgb_c_1));
    InMux I__965 (
            .O(N__12782),
            .I(N__12779));
    LocalMux I__964 (
            .O(N__12779),
            .I(\this_delay_clk.M_pipe_qZ0Z_1 ));
    InMux I__963 (
            .O(N__12776),
            .I(N__12773));
    LocalMux I__962 (
            .O(N__12773),
            .I(\this_delay_clk.M_pipe_qZ0Z_2 ));
    IoInMux I__961 (
            .O(N__12770),
            .I(N__12767));
    LocalMux I__960 (
            .O(N__12767),
            .I(N__12764));
    Odrv12 I__959 (
            .O(N__12764),
            .I(rgb_c_2));
    IoInMux I__958 (
            .O(N__12761),
            .I(N__12758));
    LocalMux I__957 (
            .O(N__12758),
            .I(N__12755));
    Span4Mux_s3_h I__956 (
            .O(N__12755),
            .I(N__12752));
    Span4Mux_v I__955 (
            .O(N__12752),
            .I(N__12749));
    Span4Mux_v I__954 (
            .O(N__12749),
            .I(N__12746));
    Odrv4 I__953 (
            .O(N__12746),
            .I(rgb_c_4));
    IoInMux I__952 (
            .O(N__12743),
            .I(N__12740));
    LocalMux I__951 (
            .O(N__12740),
            .I(N__12737));
    Span4Mux_s3_h I__950 (
            .O(N__12737),
            .I(N__12734));
    Span4Mux_v I__949 (
            .O(N__12734),
            .I(N__12731));
    Odrv4 I__948 (
            .O(N__12731),
            .I(rgb_c_5));
    CascadeMux I__947 (
            .O(N__12728),
            .I(N__12725));
    InMux I__946 (
            .O(N__12725),
            .I(N__12722));
    LocalMux I__945 (
            .O(N__12722),
            .I(N__12719));
    Odrv12 I__944 (
            .O(N__12719),
            .I(M_this_vga_signals_address_6));
    IoInMux I__943 (
            .O(N__12716),
            .I(N__12713));
    LocalMux I__942 (
            .O(N__12713),
            .I(port_data_rw_0_i));
    InMux I__941 (
            .O(N__12710),
            .I(N__12707));
    LocalMux I__940 (
            .O(N__12707),
            .I(N__12704));
    Span4Mux_v I__939 (
            .O(N__12704),
            .I(N__12701));
    Odrv4 I__938 (
            .O(N__12701),
            .I(port_clk_c));
    InMux I__937 (
            .O(N__12698),
            .I(N__12695));
    LocalMux I__936 (
            .O(N__12695),
            .I(\this_delay_clk.M_pipe_qZ0Z_0 ));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\this_ppu.un1_M_surface_y_d_cry_6 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_8),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_16),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(un1_M_this_warmup_d_cry_24),
            .carryinitout(bfn_10_23_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_15_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_20_0_ (
            .carryinitin(M_this_data_count_q_cry_7),
            .carryinitout(bfn_15_20_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_21_24_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_24_0_));
    defparam IN_MUX_bfv_21_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_25_0_ (
            .carryinitin(un1_M_this_ext_address_q_cry_7),
            .carryinitout(bfn_21_25_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(un1_M_this_spr_address_q_cry_7),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_26_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_26_25_0_));
    defparam IN_MUX_bfv_26_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_26_26_0_ (
            .carryinitin(un1_M_this_map_address_q_cry_7),
            .carryinitout(bfn_26_26_0_));
    ICE_GB \this_vga_signals.M_vcounter_q_esr_RNINK957_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__29654),
            .GLOBALBUFFEROUTPUT(\this_vga_signals.N_1188_g ));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_9  (
            .USERSIGNALTOGLOBALBUFFER(N__31013),
            .GLOBALBUFFEROUTPUT(M_this_reset_cond_out_g_0));
    ICE_GB \this_reset_cond.M_stage_q_RNIC5C7_0_9  (
            .USERSIGNALTOGLOBALBUFFER(N__30125),
            .GLOBALBUFFEROUTPUT(N_527_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.port_data_rw_0_i_LC_1_21_7 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \this_vga_signals.port_data_rw_0_i_LC_1_21_7  (
            .in0(N__34178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31540),
            .lcout(port_data_rw_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_1_LC_2_19_1 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_1_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_1_LC_2_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_1_LC_2_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12698),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39414),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_0_LC_2_19_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_0_LC_2_19_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_0_LC_2_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_delay_clk.M_pipe_q_0_LC_2_19_5  (
            .in0(N__12710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39414),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_18_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__14654),
            .in2(_gnd_net_),
            .in3(N__13776),
            .lcout(rgb_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_4  (
            .in0(N__13775),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13064),
            .lcout(rgb_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_2 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_2 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_3_LC_3_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_3_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12776),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39410),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_3 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_2_LC_3_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_2_LC_3_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12782),
            .lcout(\this_delay_clk.M_pipe_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39410),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_0  (
            .in0(N__14426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13760),
            .lcout(rgb_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_4_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_4_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_4_19_5 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_4_19_5  (
            .in0(N__15596),
            .in1(N__13868),
            .in2(N__13850),
            .in3(N__15539),
            .lcout(\this_vga_signals.un2_hsynclto6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_20_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_20_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_20_0  (
            .in0(N__13777),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14630),
            .lcout(rgb_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_21_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_21_4  (
            .in0(N__13781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14453),
            .lcout(rgb_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFI285_9_LC_5_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFI285_9_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIFI285_9_LC_5_17_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIFI285_9_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__12827),
            .in2(_gnd_net_),
            .in3(N__26468),
            .lcout(M_this_vga_signals_address_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_5_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_5_17_1 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_5_17_1  (
            .in0(N__13917),
            .in1(N__13184),
            .in2(N__13985),
            .in3(N__12959),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1 ),
            .ltout(\this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_1_LC_5_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_1_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_1_LC_5_17_2 .LUT_INIT=16'b0010010001000010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_1_LC_5_17_2  (
            .in0(N__15581),
            .in1(N__15531),
            .in2(N__12872),
            .in3(N__12859),
            .lcout(\this_vga_signals.mult1_un89_sum_c3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_0_LC_5_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_0_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_0_LC_5_17_3 .LUT_INIT=16'b1101001001001011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_0_LC_5_17_3  (
            .in0(N__13039),
            .in1(N__15582),
            .in2(N__12821),
            .in3(N__13916),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_5_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_5_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__12850),
            .in2(N__12869),
            .in3(N__12860),
            .lcout(\this_vga_signals.mult1_un89_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_LC_5_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_LC_5_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_LC_5_17_5 .LUT_INIT=16'b1100110010010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_LC_5_17_5  (
            .in0(N__13040),
            .in1(N__15583),
            .in2(N__13924),
            .in3(N__12866),
            .lcout(\this_vga_signals.mult1_un89_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_5_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_5_17_6 .LUT_INIT=16'b1001101110001001;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_5_17_6  (
            .in0(N__13915),
            .in1(N__12817),
            .in2(N__15591),
            .in3(N__13038),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un82_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNISNQ4B1_9_LC_5_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNISNQ4B1_9_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNISNQ4B1_9_LC_5_17_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNISNQ4B1_9_LC_5_17_7  (
            .in0(N__12851),
            .in1(_gnd_net_),
            .in2(N__12842),
            .in3(N__26469),
            .lcout(M_this_vga_signals_address_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_5_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_5_18_0 .LUT_INIT=16'b1101010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_5_18_0  (
            .in0(N__14173),
            .in1(N__14103),
            .in2(N__14243),
            .in3(N__14295),
            .lcout(\this_vga_signals.SUM_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_5_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_5_18_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__13973),
            .in2(_gnd_net_),
            .in3(N__13183),
            .lcout(\this_vga_signals.mult1_un75_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_2_LC_5_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_2_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_2_LC_5_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_2_LC_5_18_3  (
            .in0(N__13845),
            .in1(N__13138),
            .in2(N__13983),
            .in3(N__13037),
            .lcout(\this_vga_signals.mult1_un82_sum_axbxc3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_5_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_5_18_4 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_5_18_4  (
            .in0(N__12953),
            .in1(N__14104),
            .in2(N__14375),
            .in3(N__14296),
            .lcout(\this_vga_signals.hsync_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_5_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_5_18_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_5_18_5  (
            .in0(N__13846),
            .in1(N__15592),
            .in2(N__13984),
            .in3(N__13925),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclt7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_5_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_5_18_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_5_18_6  (
            .in0(N__14374),
            .in1(N__14105),
            .in2(N__12947),
            .in3(N__14297),
            .lcout(),
            .ltout(\this_vga_signals.un4_hsynclt8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_5_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_5_18_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_5_18_7  (
            .in0(N__12944),
            .in1(N__14240),
            .in2(N__12938),
            .in3(N__14174),
            .lcout(this_vga_signals_hsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNICT164_9_LC_5_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICT164_9_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNICT164_9_LC_5_19_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNICT164_9_LC_5_19_6  (
            .in0(N__14241),
            .in1(N__14171),
            .in2(N__29618),
            .in3(N__14101),
            .lcout(M_this_vga_ramdac_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_5_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_5_20_5 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_5_20_5  (
            .in0(N__14102),
            .in1(N__14242),
            .in2(_gnd_net_),
            .in3(N__14172),
            .lcout(this_vga_signals_hvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_0_9_LC_5_24_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_0_9_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_0_9_LC_5_24_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_0_9_LC_5_24_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29617),
            .lcout(this_vga_signals_vvisibility_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_16_0 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_16_0  (
            .in0(N__13768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14405),
            .lcout(rgb_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_17_0 .LUT_INIT=16'b1001111011010110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_17_0  (
            .in0(N__14359),
            .in1(N__12970),
            .in2(N__13844),
            .in3(N__13111),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1 .LUT_INIT=16'b0111101000011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1  (
            .in0(N__13968),
            .in1(N__13899),
            .in2(N__13043),
            .in3(N__13004),
            .lcout(\this_vga_signals.mult1_un75_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un75_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUG6BC_9_LC_6_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUG6BC_9_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIUG6BC_9_LC_6_17_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIUG6BC_9_LC_6_17_2  (
            .in0(N__26481),
            .in1(_gnd_net_),
            .in2(N__13022),
            .in3(_gnd_net_),
            .lcout(M_this_vga_signals_address_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_1_LC_6_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_1_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_1_LC_6_17_3 .LUT_INIT=16'b0101000011110101;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_1_LC_6_17_3  (
            .in0(N__13110),
            .in1(_gnd_net_),
            .in2(N__14361),
            .in3(N__13831),
            .lcout(),
            .ltout(\this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_LC_6_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_LC_6_17_4 .LUT_INIT=16'b1000010101011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_LC_6_17_4  (
            .in0(N__14276),
            .in1(N__14349),
            .in2(N__13007),
            .in3(N__13091),
            .lcout(\this_vga_signals.if_m7_0_o4_1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_6_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_6_17_5 .LUT_INIT=16'b1001010111010111;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_6_17_5  (
            .in0(N__14140),
            .in1(N__14068),
            .in2(N__14218),
            .in3(N__14274),
            .lcout(\this_vga_signals.SUM_3 ),
            .ltout(\this_vga_signals.SUM_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_17_6 .LUT_INIT=16'b0101101001011110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_17_6  (
            .in0(N__14275),
            .in1(N__14345),
            .in2(N__12998),
            .in3(N__13109),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73OIC3_9_LC_6_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73OIC3_9_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI73OIC3_9_LC_6_17_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI73OIC3_9_LC_6_17_7  (
            .in0(N__12995),
            .in1(N__26480),
            .in2(_gnd_net_),
            .in3(N__12989),
            .lcout(M_this_vga_signals_address_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_6_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_6_18_0 .LUT_INIT=16'b0110111000100110;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_6_18_0  (
            .in0(N__14358),
            .in1(N__12971),
            .in2(N__13840),
            .in3(N__13112),
            .lcout(\this_vga_signals.mult1_un61_sum_axbxc3_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_LC_6_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_LC_6_18_1 .LUT_INIT=16'b1111110101000000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_LC_6_18_1  (
            .in0(N__13959),
            .in1(N__13825),
            .in2(N__13187),
            .in3(N__13070),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_2 ),
            .ltout(\this_vga_signals.mult1_un68_sum_c3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0J6BC_9_LC_6_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0J6BC_9_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI0J6BC_9_LC_6_18_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI0J6BC_9_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13172),
            .in3(N__26460),
            .lcout(M_this_vga_signals_address_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRU9S6_9_LC_6_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRU9S6_9_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIRU9S6_9_LC_6_18_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIRU9S6_9_LC_6_18_3  (
            .in0(N__26462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13079),
            .lcout(M_this_vga_signals_address_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI59HG8_9_LC_6_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI59HG8_9_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI59HG8_9_LC_6_18_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI59HG8_9_LC_6_18_4  (
            .in0(_gnd_net_),
            .in1(N__26461),
            .in2(_gnd_net_),
            .in3(N__13139),
            .lcout(M_this_vga_signals_address_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_6_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_6_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_6_18_5 .LUT_INIT=16'b0100001010111101;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_6_18_5  (
            .in0(N__14139),
            .in1(N__14067),
            .in2(N__14217),
            .in3(N__14272),
            .lcout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9 ),
            .ltout(\this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_6 .LUT_INIT=16'b1111001010110000;
    LogicCell40 \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_6  (
            .in0(N__14273),
            .in1(N__14350),
            .in2(N__13094),
            .in3(N__13090),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un4_haddress_if_m1_1_LC_6_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un4_haddress_if_m1_1_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un4_haddress_if_m1_1_LC_6_18_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un4_haddress_if_m1_1_LC_6_18_7  (
            .in0(N__14351),
            .in1(_gnd_net_),
            .in2(N__13073),
            .in3(N__13821),
            .lcout(\this_vga_signals.if_m1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_19_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_19_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_19_2 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_19_2  (
            .in0(N__14501),
            .in1(N__31014),
            .in2(N__13060),
            .in3(N__16169),
            .lcout(\this_vga_ramdac.N_3139_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39398),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_7_17_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_7_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__15584),
            .in2(N__15538),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_17_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_2_LC_7_17_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_2_LC_7_17_1  (
            .in0(N__29783),
            .in1(N__13911),
            .in2(_gnd_net_),
            .in3(N__13211),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_1 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_17_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_3_LC_7_17_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_3_LC_7_17_2  (
            .in0(N__29787),
            .in1(N__13972),
            .in2(_gnd_net_),
            .in3(N__13208),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_2 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_17_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_4_LC_7_17_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_4_LC_7_17_3  (
            .in0(N__29784),
            .in1(N__13826),
            .in2(_gnd_net_),
            .in3(N__13205),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_3 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_17_4 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_5_LC_7_17_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_5_LC_7_17_4  (
            .in0(N__29788),
            .in1(N__14360),
            .in2(_gnd_net_),
            .in3(N__13202),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_4 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_17_5 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_6_LC_7_17_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_6_LC_7_17_5  (
            .in0(N__29785),
            .in1(N__14283),
            .in2(_gnd_net_),
            .in3(N__13199),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_6 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_5 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_7_LC_7_17_6 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_7_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_7_LC_7_17_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_7_LC_7_17_6  (
            .in0(N__29789),
            .in1(N__14077),
            .in2(_gnd_net_),
            .in3(N__13196),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_7 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_6 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_8_LC_7_17_7 .C_ON=1'b1;
    defparam \this_vga_signals.M_hcounter_q_8_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_8_LC_7_17_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_8_LC_7_17_7  (
            .in0(N__29786),
            .in1(N__14149),
            .in2(_gnd_net_),
            .in3(N__13193),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_8 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_hcounter_d_cry_7 ),
            .carryout(\this_vga_signals.un1_M_hcounter_d_cry_8 ),
            .clk(N__39381),
            .ce(),
            .sr(N__16289));
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_esr_9_LC_7_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_9_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__14216),
            .in2(_gnd_net_),
            .in3(N__13190),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39386),
            .ce(N__16259),
            .sr(N__16285));
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_7_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_e_0_LC_7_19_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_0_LC_7_19_0  (
            .in0(N__16313),
            .in1(N__16247),
            .in2(_gnd_net_),
            .in3(N__28615),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39393),
            .ce(N__29792),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_7_19_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_7_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__13334),
            .in2(_gnd_net_),
            .in3(N__23988),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_7_19_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_7_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_7_19_2  (
            .in0(N__23989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13310),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_7_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_7_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__23992),
            .in2(_gnd_net_),
            .in3(N__13541),
            .lcout(\this_ppu.oam_cache.N_823_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_7_19_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_7_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_7_19_4  (
            .in0(N__23990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13583),
            .lcout(\this_ppu.oam_cache.N_820_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_7_19_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_7_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_7_19_5  (
            .in0(N__13277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23993),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_7_19_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_7_19_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_7_19_6  (
            .in0(N__23991),
            .in1(N__13253),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_7_19_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_7_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__13232),
            .in2(_gnd_net_),
            .in3(N__23994),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_7_20_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_7_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__23987),
            .in2(N__13449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_20_0_),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_7_20_1 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(N__13359),
            .in2(_gnd_net_),
            .in3(N__13214),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_0 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_7_20_2 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_7_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13408),
            .in3(N__13484),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_1 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_7_20_3 .C_ON=1'b1;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_7_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(N__13700),
            .in2(_gnd_net_),
            .in3(N__13481),
            .lcout(\this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\this_ppu.un1_M_oam_cache_cnt_q_cry_2 ),
            .carryout(\this_ppu.un1_M_oam_cache_cnt_q_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_7_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_4_LC_7_20_4 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_4_LC_7_20_4  (
            .in0(N__13475),
            .in1(N__21623),
            .in2(N__21524),
            .in3(N__13478),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39399),
            .ce(),
            .sr(N__38962));
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_1_LC_7_21_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_1_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_1_LC_7_21_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m71_i_o2_1_LC_7_21_0  (
            .in0(N__13358),
            .in1(N__18247),
            .in2(N__13704),
            .in3(N__18407),
            .lcout(\this_ppu.m71_i_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_0_LC_7_21_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_0_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_0_LC_7_21_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m71_i_o2_0_LC_7_21_1  (
            .in0(N__13442),
            .in1(N__18339),
            .in2(N__13407),
            .in3(N__18544),
            .lcout(),
            .ltout(\this_ppu.m71_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_LC_7_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_o2_LC_7_21_2 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m71_i_o2_LC_7_21_2  (
            .in0(N__18670),
            .in1(N__13474),
            .in2(N__13463),
            .in3(N__13460),
            .lcout(\this_ppu.N_796_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_7_21_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_0_LC_7_21_3 .LUT_INIT=16'b0001001001011010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_0_LC_7_21_3  (
            .in0(N__23983),
            .in1(N__21612),
            .in2(N__13450),
            .in3(N__21522),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39404),
            .ce(),
            .sr(N__38959));
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_7_21_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_2_LC_7_21_4 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_2_LC_7_21_4  (
            .in0(N__21520),
            .in1(N__13418),
            .in2(N__21622),
            .in3(N__13400),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39404),
            .ce(),
            .sr(N__38959));
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_7_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_1_LC_7_21_5 .LUT_INIT=16'b0001001001011010;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_1_LC_7_21_5  (
            .in0(N__13360),
            .in1(N__21613),
            .in2(N__13376),
            .in3(N__21523),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39404),
            .ce(),
            .sr(N__38959));
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_7_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_cache_cnt_q_3_LC_7_21_6 .LUT_INIT=16'b0001010000111100;
    LogicCell40 \this_ppu.M_oam_cache_cnt_q_3_LC_7_21_6  (
            .in0(N__21521),
            .in1(N__13715),
            .in2(N__13705),
            .in3(N__21620),
            .lcout(\this_ppu.M_oam_cache_cnt_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39404),
            .ce(),
            .sr(N__38959));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_7_21_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_7_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_7_21_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_7_21_7  (
            .in0(N__23982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13604),
            .lcout(\this_ppu.oam_cache.N_826_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_24_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_24_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_24_3  (
            .in0(_gnd_net_),
            .in1(N__23978),
            .in2(_gnd_net_),
            .in3(N__14018),
            .lcout(\this_ppu.oam_cache.N_824_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_7_24_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_7_24_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_7_24_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_7_24_4  (
            .in0(N__23981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14036),
            .lcout(\this_ppu.oam_cache.N_821_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_7_24_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_7_24_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_7_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_7_24_5  (
            .in0(_gnd_net_),
            .in1(N__23979),
            .in2(_gnd_net_),
            .in3(N__13502),
            .lcout(\this_ppu.oam_cache.N_822_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_24_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_24_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_24_6  (
            .in0(N__23980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13520),
            .lcout(\this_ppu.oam_cache.N_819_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_7_24_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_7_24_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_7_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_7_24_7  (
            .in0(_gnd_net_),
            .in1(N__23977),
            .in2(_gnd_net_),
            .in3(N__13562),
            .lcout(\this_ppu.oam_cache.N_825_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_4_LC_7_28_2 .C_ON=1'b0;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_4_LC_7_28_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_4_LC_7_28_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.un1_M_state_q_7_i_a2_7_4_LC_7_28_2  (
            .in0(N__13597),
            .in1(N__13579),
            .in2(N__13561),
            .in3(N__13534),
            .lcout(\this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_3_LC_7_28_5 .C_ON=1'b0;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_3_LC_7_28_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_3_LC_7_28_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_ppu.un1_M_state_q_7_i_a2_7_3_LC_7_28_5  (
            .in0(_gnd_net_),
            .in1(N__13516),
            .in2(_gnd_net_),
            .in3(N__13498),
            .lcout(),
            .ltout(\this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_LC_7_28_6 .C_ON=1'b0;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_state_q_7_i_a2_7_LC_7_28_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.un1_M_state_q_7_i_a2_7_LC_7_28_6  (
            .in0(N__14032),
            .in1(N__14014),
            .in2(N__14000),
            .in3(N__13997),
            .lcout(\this_ppu.N_838_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_a2_0_LC_9_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_a2_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m48_i_a2_0_LC_9_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m48_i_a2_0_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__24050),
            .in2(_gnd_net_),
            .in3(N__21784),
            .lcout(\this_ppu.m48_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_11_LC_9_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_11_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_11_LC_9_16_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.M_state_q_11_LC_9_16_0  (
            .in0(N__21377),
            .in1(N__21722),
            .in2(_gnd_net_),
            .in3(N__36959),
            .lcout(\this_ppu.M_state_qZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39357),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_3_LC_9_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_3_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_3_LC_9_16_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_a2_3_LC_9_16_2  (
            .in0(N__17089),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18860),
            .lcout(),
            .ltout(\this_ppu.m35_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_LC_9_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_LC_9_16_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_a2_LC_9_16_3  (
            .in0(N__18240),
            .in1(N__18666),
            .in2(N__13991),
            .in3(N__16814),
            .lcout(\this_ppu.N_802 ),
            .ltout(\this_ppu.N_802_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_2_LC_9_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_2_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_2_LC_9_16_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \this_ppu.M_state_q_2_LC_9_16_4  (
            .in0(N__17090),
            .in1(_gnd_net_),
            .in2(N__13988),
            .in3(N__36960),
            .lcout(\this_ppu.M_state_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39357),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_9_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_9_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_9_17_0  (
            .in0(_gnd_net_),
            .in1(N__13960),
            .in2(_gnd_net_),
            .in3(N__13900),
            .lcout(\this_vga_signals.un2_hsynclto3_1 ),
            .ltout(\this_vga_signals.un2_hsynclto3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_9_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_9_17_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_9_17_1  (
            .in0(N__15559),
            .in1(N__15519),
            .in2(N__13853),
            .in3(N__13830),
            .lcout(\this_vga_signals.M_hcounter_d7lt7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_17_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_q_ret_LC_9_17_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_q_ret_LC_9_17_2  (
            .in0(N__30985),
            .in1(N__26491),
            .in2(N__13767),
            .in3(N__16159),
            .lcout(\this_vga_ramdac.M_this_vga_ramdac_en_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39366),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_17_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_17_3 .LUT_INIT=16'b0001010100101111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_17_3  (
            .in0(N__14530),
            .in1(N__14609),
            .in2(N__14585),
            .in3(N__14560),
            .lcout(),
            .ltout(\this_vga_ramdac.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_17_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_17_4 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_17_4  (
            .in0(N__30987),
            .in1(N__14422),
            .in2(N__14429),
            .in3(N__16158),
            .lcout(\this_vga_ramdac.N_3140_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39366),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_17_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_17_5 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_17_5  (
            .in0(N__14531),
            .in1(N__14559),
            .in2(_gnd_net_),
            .in3(N__14608),
            .lcout(),
            .ltout(\this_vga_ramdac.N_24_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_17_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_17_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_17_6  (
            .in0(N__30986),
            .in1(N__14398),
            .in2(N__14408),
            .in3(N__16157),
            .lcout(\this_vga_ramdac.N_3138_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39366),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_6_LC_9_17_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_6_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_6_LC_9_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_6_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14387),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39366),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIVCD62_9_LC_9_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIVCD62_9_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIVCD62_9_LC_9_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIVCD62_9_LC_9_18_0  (
            .in0(N__14370),
            .in1(N__14219),
            .in2(N__14306),
            .in3(N__14294),
            .lcout(),
            .ltout(\this_vga_signals.N_864_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNITLAV2_9_LC_9_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNITLAV2_9_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNITLAV2_9_LC_9_18_1 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNITLAV2_9_LC_9_18_1  (
            .in0(N__14220),
            .in1(N__14165),
            .in2(N__14108),
            .in3(N__14093),
            .lcout(\this_vga_signals.M_hcounter_d7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_18_2 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_18_2 .LUT_INIT=16'b0000101110010111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_18_2  (
            .in0(N__14580),
            .in1(N__14557),
            .in2(N__14533),
            .in3(N__14606),
            .lcout(),
            .ltout(\this_vga_ramdac.m16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_18_3 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_18_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_18_3  (
            .in0(N__14644),
            .in1(N__30988),
            .in2(N__14657),
            .in3(N__16164),
            .lcout(\this_vga_ramdac.N_3141_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39374),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_18_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_18_4 .LUT_INIT=16'b0101100100101011;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_18_4  (
            .in0(N__14581),
            .in1(N__14558),
            .in2(N__14534),
            .in3(N__14607),
            .lcout(),
            .ltout(\this_vga_ramdac.m19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_5 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_5 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_5  (
            .in0(N__14620),
            .in1(N__30989),
            .in2(N__14633),
            .in3(N__16165),
            .lcout(\this_vga_ramdac.N_3142_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39374),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_6 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_6 .LUT_INIT=16'b0101001100011001;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_6  (
            .in0(N__14579),
            .in1(N__14556),
            .in2(N__14532),
            .in3(N__14605),
            .lcout(\this_vga_ramdac.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_18_7 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_18_7 .LUT_INIT=16'b0011001000111111;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_18_7  (
            .in0(N__14604),
            .in1(N__14578),
            .in2(N__14561),
            .in3(N__14520),
            .lcout(\this_vga_ramdac.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_9_19_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNID8M7_17_LC_9_19_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNID8M7_17_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14477),
            .lcout(\this_ppu.M_oam_cache_read_data_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_17_LC_9_19_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_17_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_17_LC_9_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_17_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14489),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39382),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_16_LC_9_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_16_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_16_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_16_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14471),
            .lcout(\this_ppu.M_oam_cache_read_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39382),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_19_4 .C_ON=1'b0;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_19_4 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_19_4  (
            .in0(N__14459),
            .in1(N__30991),
            .in2(N__14446),
            .in3(N__16160),
            .lcout(\this_vga_ramdac.N_3143_reto ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39382),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_9_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_0_1_LC_9_19_5 .LUT_INIT=16'b0010001001100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_1_LC_9_19_5  (
            .in0(N__16243),
            .in1(N__29774),
            .in2(N__16219),
            .in3(N__28586),
            .lcout(\this_vga_signals.M_pcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39382),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_18_LC_9_19_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_18_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_18_LC_9_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_18_LC_9_19_7  (
            .in0(N__14744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39382),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIC31GS_2_LC_9_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIC31GS_2_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIC31GS_2_LC_9_20_0 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIC31GS_2_LC_9_20_0  (
            .in0(N__18408),
            .in1(N__18800),
            .in2(N__18350),
            .in3(N__18452),
            .lcout(\this_ppu.N_777_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIKRNBS_1_LC_9_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIKRNBS_1_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIKRNBS_1_LC_9_20_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIKRNBS_1_LC_9_20_2  (
            .in0(N__18409),
            .in1(N__18798),
            .in2(_gnd_net_),
            .in3(N__18451),
            .lcout(\this_ppu.N_776_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_LC_9_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_LC_9_20_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_LC_9_20_3  (
            .in0(N__14774),
            .in1(N__14762),
            .in2(N__14786),
            .in3(N__14804),
            .lcout(\this_ppu.N_932_0 ),
            .ltout(\this_ppu.N_932_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_0_LC_9_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_0_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_0_LC_9_20_4 .LUT_INIT=16'b0001000100110001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_0_LC_9_20_4  (
            .in0(N__17258),
            .in1(N__23849),
            .in2(N__14705),
            .in3(N__14677),
            .lcout(\this_ppu.un1_M_state_q_7_i_0_0 ),
            .ltout(\this_ppu.un1_M_state_q_7_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNITKE7S_0_LC_9_20_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNITKE7S_0_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNITKE7S_0_LC_9_20_5 .LUT_INIT=16'b1000001000100010;
    LogicCell40 \this_ppu.M_oam_curr_q_RNITKE7S_0_LC_9_20_5  (
            .in0(N__18799),
            .in1(N__18540),
            .in2(N__14702),
            .in3(N__18578),
            .lcout(\this_ppu.N_775_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_3_LC_9_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_3_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_3_LC_9_20_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_3_LC_9_20_6  (
            .in0(N__17259),
            .in1(N__14684),
            .in2(_gnd_net_),
            .in3(N__14678),
            .lcout(\this_ppu.M_state_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39389),
            .ce(),
            .sr(N__36831));
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_9_21_0 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_9_21_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__14663),
            .in2(N__22742),
            .in3(N__23482),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\this_ppu.un1_oam_data_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_9_21_1 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_9_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__14816),
            .in2(N__22694),
            .in3(N__23437),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_17 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_0 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_9_21_2 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_9_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__14810),
            .in2(N__22652),
            .in3(N__23398),
            .lcout(\this_ppu.M_this_oam_ram_read_data_i_18 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_1 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_0_LC_9_21_3 .C_ON=1'b1;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_0_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_0_LC_9_21_3 .LUT_INIT=16'b0001010001000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_0_LC_9_21_3  (
            .in0(N__14795),
            .in1(N__15116),
            .in2(N__22606),
            .in3(N__14798),
            .lcout(\this_ppu.m28_e_i_o2_0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_2 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_9_21_4 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__15482),
            .in2(N__22555),
            .in3(N__14789),
            .lcout(\this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_3 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_9_21_5 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__14996),
            .in2(N__22495),
            .in3(N__14777),
            .lcout(\this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_4 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_9_21_6 .C_ON=1'b1;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__14954),
            .in2(N__22438),
            .in3(N__14768),
            .lcout(\this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0 ),
            .ltout(),
            .carryin(\this_ppu.un1_oam_data_1_cry_5 ),
            .carryout(\this_ppu.un1_oam_data_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLD_LC_9_21_7 .C_ON=1'b0;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLD_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLD_LC_9_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLD_LC_9_21_7  (
            .in0(N__14947),
            .in1(N__23296),
            .in2(_gnd_net_),
            .in3(N__14765),
            .lcout(\this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_22_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_22_0  (
            .in0(N__23884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15017),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_22_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_22_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_22_2  (
            .in0(N__14972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23885),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_22_3 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_22_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14971),
            .lcout(M_this_oam_ram_read_data_i_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_9_22_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_9_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__23886),
            .in2(_gnd_net_),
            .in3(N__14948),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_9_22_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_9_22_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(N__23883),
            .in2(_gnd_net_),
            .in3(N__14918),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_22_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_22_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(N__14891),
            .in2(_gnd_net_),
            .in3(N__23887),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_9_22_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_9_22_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_9_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(N__23882),
            .in2(_gnd_net_),
            .in3(N__14870),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_6_LC_9_27_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_6_LC_9_27_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_6_LC_9_27_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_6_LC_9_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37389),
            .lcout(M_this_data_tmp_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39420),
            .ce(N__23620),
            .sr(N__36841));
    defparam M_this_data_tmp_q_esr_3_LC_9_27_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_3_LC_9_27_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_3_LC_9_27_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_3_LC_9_27_7 (
            .in0(N__37860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39420),
            .ce(N__23620),
            .sr(N__36841));
    defparam \this_start_data_delay.M_last_q_RNIPR151_LC_9_28_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIPR151_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIPR151_LC_9_28_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIPR151_LC_9_28_0  (
            .in0(N__19370),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16661),
            .lcout(M_this_oam_ram_write_data_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_9_28_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_9_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_9_28_1  (
            .in0(_gnd_net_),
            .in1(N__14840),
            .in2(_gnd_net_),
            .in3(N__23972),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOQ151_LC_9_28_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOQ151_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOQ151_LC_9_28_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOQ151_LC_9_28_3  (
            .in0(_gnd_net_),
            .in1(N__17153),
            .in2(_gnd_net_),
            .in3(N__19373),
            .lcout(M_this_oam_ram_write_data_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIQS151_LC_9_28_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIQS151_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIQS151_LC_9_28_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIQS151_LC_9_28_4  (
            .in0(N__19371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17162),
            .lcout(M_this_oam_ram_write_data_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNITV151_LC_9_28_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNITV151_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNITV151_LC_9_28_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNITV151_LC_9_28_5  (
            .in0(_gnd_net_),
            .in1(N__21881),
            .in2(_gnd_net_),
            .in3(N__19369),
            .lcout(M_this_oam_ram_write_data_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_9_28_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_9_28_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_9_28_6  (
            .in0(N__23971),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15062),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICRDD1_LC_9_28_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICRDD1_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICRDD1_LC_9_28_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNICRDD1_LC_9_28_7  (
            .in0(_gnd_net_),
            .in1(N__16667),
            .in2(_gnd_net_),
            .in3(N__19372),
            .lcout(M_this_oam_ram_write_data_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI7MDD1_LC_9_29_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI7MDD1_LC_9_29_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI7MDD1_LC_9_29_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI7MDD1_LC_9_29_0  (
            .in0(N__19375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15032),
            .lcout(M_this_oam_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_9_29_1 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_9_29_1 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_9_29_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_9_29_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15013),
            .lcout(M_this_oam_ram_read_data_i_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIAPDD1_LC_9_29_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIAPDD1_LC_9_29_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIAPDD1_LC_9_29_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIAPDD1_LC_9_29_2  (
            .in0(N__19377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14987),
            .lcout(M_this_oam_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI9ODD1_LC_9_29_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI9ODD1_LC_9_29_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI9ODD1_LC_9_29_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI9ODD1_LC_9_29_4  (
            .in0(N__19376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16619),
            .lcout(M_this_oam_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBQDD1_LC_9_29_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBQDD1_LC_9_29_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBQDD1_LC_9_29_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBQDD1_LC_9_29_5  (
            .in0(_gnd_net_),
            .in1(N__16625),
            .in2(_gnd_net_),
            .in3(N__19374),
            .lcout(M_this_oam_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_9_30_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_9_30_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_9_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_9_30_0  (
            .in0(_gnd_net_),
            .in1(N__15197),
            .in2(_gnd_net_),
            .in3(N__23973),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_9_30_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_9_30_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_9_30_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_9_30_1  (
            .in0(N__23975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15176),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIRT151_LC_9_30_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIRT151_LC_9_30_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIRT151_LC_9_30_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIRT151_LC_9_30_2  (
            .in0(_gnd_net_),
            .in1(N__19365),
            .in2(_gnd_net_),
            .in3(N__16607),
            .lcout(M_this_oam_ram_write_data_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOR251_LC_9_30_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOR251_LC_9_30_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOR251_LC_9_30_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOR251_LC_9_30_3  (
            .in0(N__16613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19378),
            .lcout(M_this_oam_ram_write_data_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_9_30_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_9_30_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_9_30_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_9_30_4  (
            .in0(N__15128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23976),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_30_5 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_30_5 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_30_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_30_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15127),
            .lcout(M_this_oam_ram_read_data_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_9_30_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_9_30_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_9_30_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_9_30_6  (
            .in0(N__15494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23974),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_30_7 .C_ON=1'b0;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_30_7 .SEQ_MODE=4'b0000;
    defparam \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_30_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_30_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15493),
            .lcout(M_this_oam_ram_read_data_i_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI43IG1_LC_9_31_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI43IG1_LC_9_31_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI43IG1_LC_9_31_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI43IG1_LC_9_31_0  (
            .in0(N__19380),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37853),
            .lcout(M_this_oam_ram_write_data_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI76IG1_LC_9_31_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI76IG1_LC_9_31_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI76IG1_LC_9_31_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI76IG1_LC_9_31_3  (
            .in0(_gnd_net_),
            .in1(N__37397),
            .in2(_gnd_net_),
            .in3(N__19382),
            .lcout(M_this_oam_ram_write_data_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNISU151_LC_9_31_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNISU151_LC_9_31_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNISU151_LC_9_31_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNISU151_LC_9_31_4  (
            .in0(N__19383),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17540),
            .lcout(M_this_oam_ram_write_data_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI65IG1_LC_9_31_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI65IG1_LC_9_31_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI65IG1_LC_9_31_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI65IG1_LC_9_31_5  (
            .in0(N__38895),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19381),
            .lcout(M_this_oam_ram_write_data_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI10IG1_LC_9_31_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI10IG1_LC_9_31_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI10IG1_LC_9_31_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI10IG1_LC_9_31_7  (
            .in0(N__38102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19379),
            .lcout(M_this_oam_ram_write_data_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dma_0_sbtinv_LC_10_7_3.C_ON=1'b0;
    defparam dma_0_sbtinv_LC_10_7_3.SEQ_MODE=4'b0000;
    defparam dma_0_sbtinv_LC_10_7_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 dma_0_sbtinv_LC_10_7_3 (
            .in0(N__34173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dma_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_7_LC_10_10_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_7_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_7_LC_10_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_7_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15239),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39300),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_3_LC_10_12_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_3_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_3_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_3_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15224),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39309),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_4_LC_10_14_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_4_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_4_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_4_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15635),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39323),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_1_LC_10_15_1 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_1_LC_10_15_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_pixel_clk.M_counter_q_1_LC_10_15_1  (
            .in0(N__15620),
            .in1(N__15610),
            .in2(_gnd_net_),
            .in3(N__36928),
            .lcout(this_pixel_clk_M_counter_q_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39331),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.G_424_LC_10_15_5 .C_ON=1'b0;
    defparam \this_vga_signals.G_424_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.G_424_LC_10_15_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_vga_signals.G_424_LC_10_15_5  (
            .in0(N__15619),
            .in1(N__15609),
            .in2(_gnd_net_),
            .in3(N__36927),
            .lcout(\this_vga_signals.GZ0Z_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_pixel_clk.M_counter_q_0_LC_10_16_3 .C_ON=1'b0;
    defparam \this_pixel_clk.M_counter_q_0_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \this_pixel_clk.M_counter_q_0_LC_10_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_pixel_clk.M_counter_q_0_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15611),
            .lcout(this_pixel_clk_M_counter_q_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39339),
            .ce(),
            .sr(N__36825));
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_1_LC_10_17_1 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_1_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(N__15529),
            .in2(N__29779),
            .in3(N__15577),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39350),
            .ce(),
            .sr(N__16278));
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_hcounter_q_0_LC_10_17_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \this_vga_signals.M_hcounter_q_0_LC_10_17_2  (
            .in0(N__15530),
            .in1(N__29743),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_hcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39350),
            .ce(),
            .sr(N__16278));
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_17_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16364),
            .lcout(\this_ppu.M_oam_cache_read_data_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_e_RNICJLB4_0_LC_10_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNICJLB4_0_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_e_RNICJLB4_0_LC_10_18_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_e_RNICJLB4_0_LC_10_18_0  (
            .in0(N__16215),
            .in1(N__29731),
            .in2(_gnd_net_),
            .in3(N__16295),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_2_LC_10_18_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_2_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15497),
            .in3(N__16193),
            .lcout(M_this_vga_signals_pixel_clk_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39358),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_pcounter_q_ret_LC_10_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_LC_10_18_2  (
            .in0(N__16178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_pcounter_q_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39358),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_ret_RNITMRI3_LC_10_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_ret_RNITMRI3_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_ret_RNITMRI3_LC_10_18_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_vga_signals.M_pcounter_q_ret_RNITMRI3_LC_10_18_3  (
            .in0(N__16306),
            .in1(N__16241),
            .in2(_gnd_net_),
            .in3(N__28567),
            .lcout(\this_vga_signals.M_pcounter_q_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIG783_9_LC_10_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIG783_9_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNIIG783_9_LC_10_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNIIG783_9_LC_10_18_4  (
            .in0(N__28569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29732),
            .lcout(\this_vga_signals.N_1188_1 ),
            .ltout(\this_vga_signals.N_1188_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_18_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_18_5  (
            .in0(N__29734),
            .in1(_gnd_net_),
            .in2(N__16262),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.N_933_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_pcounter_q_0_RNI38654_1_LC_10_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_pcounter_q_0_RNI38654_1_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_pcounter_q_0_RNI38654_1_LC_10_18_6 .LUT_INIT=16'b0001000011001100;
    LogicCell40 \this_vga_signals.M_pcounter_q_0_RNI38654_1_LC_10_18_6  (
            .in0(N__28568),
            .in1(N__16242),
            .in2(N__16220),
            .in3(N__29733),
            .lcout(N_2_0),
            .ltout(N_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__G_462_LC_10_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__G_462_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__G_462_LC_10_18_7 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__G_462_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__16187),
            .in2(N__16181),
            .in3(N__16177),
            .lcout(G_462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_10_19_0 .C_ON=1'b1;
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_y_cry_0_c_inv_LC_10_19_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_ppu.offset_y_cry_0_c_inv_LC_10_19_0  (
            .in0(N__17512),
            .in1(N__22741),
            .in2(N__16127),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_oam_cache_read_data_i_16 ),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\this_ppu.offset_y_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_10_19_1 .C_ON=1'b1;
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_10_19_1 .LUT_INIT=16'b1100100110011100;
    LogicCell40 \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_10_19_1  (
            .in0(N__32689),
            .in1(N__22693),
            .in2(N__16118),
            .in3(N__15905),
            .lcout(M_this_ppu_spr_addr_4),
            .ltout(),
            .carryin(\this_ppu.offset_y_cry_0 ),
            .carryout(\this_ppu.offset_y_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_10_19_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_10_19_2 .LUT_INIT=16'b1100011011001001;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_10_19_2  (
            .in0(N__15902),
            .in1(N__22651),
            .in2(N__32705),
            .in3(N__15896),
            .lcout(M_this_ppu_spr_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_10_LC_10_19_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_10_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_10_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_10_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16373),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39367),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_m2_LC_10_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_m2_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m18_i_m2_LC_10_19_4 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m18_i_m2_LC_10_19_4  (
            .in0(N__17263),
            .in1(N__21568),
            .in2(N__18841),
            .in3(N__21505),
            .lcout(),
            .ltout(\this_ppu.N_836_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_1_LC_10_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_1_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_1_LC_10_19_5 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \this_ppu.M_state_q_1_LC_10_19_5  (
            .in0(N__31012),
            .in1(_gnd_net_),
            .in2(N__16355),
            .in3(N__18468),
            .lcout(\this_ppu.M_state_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39367),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_0_0_LC_10_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_0_0_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_0_0_LC_10_19_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m13_0_a2_0_0_LC_10_19_6  (
            .in0(N__21785),
            .in1(N__21721),
            .in2(_gnd_net_),
            .in3(N__21567),
            .lcout(\this_ppu.m13_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_9_LC_10_19_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_9_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_9_LC_10_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_9_LC_10_19_7  (
            .in0(N__16352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39367),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_M_this_warmup_d_cry_1_c_LC_10_20_0.C_ON=1'b1;
    defparam un1_M_this_warmup_d_cry_1_c_LC_10_20_0.SEQ_MODE=4'b0000;
    defparam un1_M_this_warmup_d_cry_1_c_LC_10_20_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_M_this_warmup_d_cry_1_c_LC_10_20_0 (
            .in0(_gnd_net_),
            .in1(N__17071),
            .in2(N__17060),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(un1_M_this_warmup_d_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_warmup_q_2_LC_10_20_1.C_ON=1'b1;
    defparam M_this_warmup_q_2_LC_10_20_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_2_LC_10_20_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_2_LC_10_20_1 (
            .in0(_gnd_net_),
            .in1(N__16340),
            .in2(_gnd_net_),
            .in3(N__16334),
            .lcout(M_this_warmup_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_1),
            .carryout(un1_M_this_warmup_d_cry_2),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_3_LC_10_20_2.C_ON=1'b1;
    defparam M_this_warmup_q_3_LC_10_20_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_3_LC_10_20_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_3_LC_10_20_2 (
            .in0(_gnd_net_),
            .in1(N__16331),
            .in2(_gnd_net_),
            .in3(N__16325),
            .lcout(M_this_warmup_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_2),
            .carryout(un1_M_this_warmup_d_cry_3),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_4_LC_10_20_3.C_ON=1'b1;
    defparam M_this_warmup_q_4_LC_10_20_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_4_LC_10_20_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_4_LC_10_20_3 (
            .in0(_gnd_net_),
            .in1(N__16322),
            .in2(_gnd_net_),
            .in3(N__16316),
            .lcout(M_this_warmup_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_3),
            .carryout(un1_M_this_warmup_d_cry_4),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_5_LC_10_20_4.C_ON=1'b1;
    defparam M_this_warmup_q_5_LC_10_20_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_5_LC_10_20_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_5_LC_10_20_4 (
            .in0(_gnd_net_),
            .in1(N__16451),
            .in2(_gnd_net_),
            .in3(N__16445),
            .lcout(M_this_warmup_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_4),
            .carryout(un1_M_this_warmup_d_cry_5),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_6_LC_10_20_5.C_ON=1'b1;
    defparam M_this_warmup_q_6_LC_10_20_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_6_LC_10_20_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_6_LC_10_20_5 (
            .in0(_gnd_net_),
            .in1(N__16442),
            .in2(_gnd_net_),
            .in3(N__16436),
            .lcout(M_this_warmup_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_5),
            .carryout(un1_M_this_warmup_d_cry_6),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_7_LC_10_20_6.C_ON=1'b1;
    defparam M_this_warmup_q_7_LC_10_20_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_7_LC_10_20_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_7_LC_10_20_6 (
            .in0(_gnd_net_),
            .in1(N__16433),
            .in2(_gnd_net_),
            .in3(N__16427),
            .lcout(M_this_warmup_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_6),
            .carryout(un1_M_this_warmup_d_cry_7),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_8_LC_10_20_7.C_ON=1'b1;
    defparam M_this_warmup_q_8_LC_10_20_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_8_LC_10_20_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_8_LC_10_20_7 (
            .in0(_gnd_net_),
            .in1(N__16424),
            .in2(_gnd_net_),
            .in3(N__16418),
            .lcout(M_this_warmup_qZ0Z_8),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_7),
            .carryout(un1_M_this_warmup_d_cry_8),
            .clk(N__39375),
            .ce(),
            .sr(N__36829));
    defparam M_this_warmup_q_9_LC_10_21_0.C_ON=1'b1;
    defparam M_this_warmup_q_9_LC_10_21_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_9_LC_10_21_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_9_LC_10_21_0 (
            .in0(_gnd_net_),
            .in1(N__16415),
            .in2(_gnd_net_),
            .in3(N__16409),
            .lcout(M_this_warmup_qZ0Z_9),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(un1_M_this_warmup_d_cry_9),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_10_LC_10_21_1.C_ON=1'b1;
    defparam M_this_warmup_q_10_LC_10_21_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_10_LC_10_21_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_10_LC_10_21_1 (
            .in0(_gnd_net_),
            .in1(N__16406),
            .in2(_gnd_net_),
            .in3(N__16400),
            .lcout(M_this_warmup_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_9),
            .carryout(un1_M_this_warmup_d_cry_10),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_11_LC_10_21_2.C_ON=1'b1;
    defparam M_this_warmup_q_11_LC_10_21_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_11_LC_10_21_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_11_LC_10_21_2 (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(_gnd_net_),
            .in3(N__16391),
            .lcout(M_this_warmup_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_10),
            .carryout(un1_M_this_warmup_d_cry_11),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_12_LC_10_21_3.C_ON=1'b1;
    defparam M_this_warmup_q_12_LC_10_21_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_12_LC_10_21_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_12_LC_10_21_3 (
            .in0(_gnd_net_),
            .in1(N__16388),
            .in2(_gnd_net_),
            .in3(N__16382),
            .lcout(M_this_warmup_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_11),
            .carryout(un1_M_this_warmup_d_cry_12),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_13_LC_10_21_4.C_ON=1'b1;
    defparam M_this_warmup_q_13_LC_10_21_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_13_LC_10_21_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_13_LC_10_21_4 (
            .in0(_gnd_net_),
            .in1(N__16379),
            .in2(_gnd_net_),
            .in3(N__16526),
            .lcout(M_this_warmup_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_12),
            .carryout(un1_M_this_warmup_d_cry_13),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_14_LC_10_21_5.C_ON=1'b1;
    defparam M_this_warmup_q_14_LC_10_21_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_14_LC_10_21_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_14_LC_10_21_5 (
            .in0(_gnd_net_),
            .in1(N__16523),
            .in2(_gnd_net_),
            .in3(N__16517),
            .lcout(M_this_warmup_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_13),
            .carryout(un1_M_this_warmup_d_cry_14),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_15_LC_10_21_6.C_ON=1'b1;
    defparam M_this_warmup_q_15_LC_10_21_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_15_LC_10_21_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_15_LC_10_21_6 (
            .in0(_gnd_net_),
            .in1(N__16514),
            .in2(_gnd_net_),
            .in3(N__16508),
            .lcout(M_this_warmup_qZ0Z_15),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_14),
            .carryout(un1_M_this_warmup_d_cry_15),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_16_LC_10_21_7.C_ON=1'b1;
    defparam M_this_warmup_q_16_LC_10_21_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_16_LC_10_21_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_16_LC_10_21_7 (
            .in0(_gnd_net_),
            .in1(N__16505),
            .in2(_gnd_net_),
            .in3(N__16499),
            .lcout(M_this_warmup_qZ0Z_16),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_15),
            .carryout(un1_M_this_warmup_d_cry_16),
            .clk(N__39383),
            .ce(),
            .sr(N__36830));
    defparam M_this_warmup_q_17_LC_10_22_0.C_ON=1'b1;
    defparam M_this_warmup_q_17_LC_10_22_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_17_LC_10_22_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_17_LC_10_22_0 (
            .in0(_gnd_net_),
            .in1(N__16496),
            .in2(_gnd_net_),
            .in3(N__16490),
            .lcout(M_this_warmup_qZ0Z_17),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(un1_M_this_warmup_d_cry_17),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_18_LC_10_22_1.C_ON=1'b1;
    defparam M_this_warmup_q_18_LC_10_22_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_18_LC_10_22_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_18_LC_10_22_1 (
            .in0(_gnd_net_),
            .in1(N__16487),
            .in2(_gnd_net_),
            .in3(N__16481),
            .lcout(M_this_warmup_qZ0Z_18),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_17),
            .carryout(un1_M_this_warmup_d_cry_18),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_19_LC_10_22_2.C_ON=1'b1;
    defparam M_this_warmup_q_19_LC_10_22_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_19_LC_10_22_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_19_LC_10_22_2 (
            .in0(_gnd_net_),
            .in1(N__16478),
            .in2(_gnd_net_),
            .in3(N__16472),
            .lcout(M_this_warmup_qZ0Z_19),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_18),
            .carryout(un1_M_this_warmup_d_cry_19),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_20_LC_10_22_3.C_ON=1'b1;
    defparam M_this_warmup_q_20_LC_10_22_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_20_LC_10_22_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_20_LC_10_22_3 (
            .in0(_gnd_net_),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__16463),
            .lcout(M_this_warmup_qZ0Z_20),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_19),
            .carryout(un1_M_this_warmup_d_cry_20),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_21_LC_10_22_4.C_ON=1'b1;
    defparam M_this_warmup_q_21_LC_10_22_4.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_21_LC_10_22_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_21_LC_10_22_4 (
            .in0(_gnd_net_),
            .in1(N__16460),
            .in2(_gnd_net_),
            .in3(N__16454),
            .lcout(M_this_warmup_qZ0Z_21),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_20),
            .carryout(un1_M_this_warmup_d_cry_21),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_22_LC_10_22_5.C_ON=1'b1;
    defparam M_this_warmup_q_22_LC_10_22_5.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_22_LC_10_22_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_22_LC_10_22_5 (
            .in0(_gnd_net_),
            .in1(N__16592),
            .in2(_gnd_net_),
            .in3(N__16586),
            .lcout(M_this_warmup_qZ0Z_22),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_21),
            .carryout(un1_M_this_warmup_d_cry_22),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_23_LC_10_22_6.C_ON=1'b1;
    defparam M_this_warmup_q_23_LC_10_22_6.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_23_LC_10_22_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_23_LC_10_22_6 (
            .in0(_gnd_net_),
            .in1(N__16583),
            .in2(_gnd_net_),
            .in3(N__16577),
            .lcout(M_this_warmup_qZ0Z_23),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_22),
            .carryout(un1_M_this_warmup_d_cry_23),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_24_LC_10_22_7.C_ON=1'b1;
    defparam M_this_warmup_q_24_LC_10_22_7.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_24_LC_10_22_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_24_LC_10_22_7 (
            .in0(_gnd_net_),
            .in1(N__16574),
            .in2(_gnd_net_),
            .in3(N__16568),
            .lcout(M_this_warmup_qZ0Z_24),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_23),
            .carryout(un1_M_this_warmup_d_cry_24),
            .clk(N__39390),
            .ce(),
            .sr(N__36832));
    defparam M_this_warmup_q_25_LC_10_23_0.C_ON=1'b1;
    defparam M_this_warmup_q_25_LC_10_23_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_25_LC_10_23_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_25_LC_10_23_0 (
            .in0(_gnd_net_),
            .in1(N__16565),
            .in2(_gnd_net_),
            .in3(N__16559),
            .lcout(M_this_warmup_qZ0Z_25),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(un1_M_this_warmup_d_cry_25),
            .clk(N__39394),
            .ce(),
            .sr(N__36833));
    defparam M_this_warmup_q_26_LC_10_23_1.C_ON=1'b1;
    defparam M_this_warmup_q_26_LC_10_23_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_26_LC_10_23_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_26_LC_10_23_1 (
            .in0(_gnd_net_),
            .in1(N__16556),
            .in2(_gnd_net_),
            .in3(N__16550),
            .lcout(M_this_warmup_qZ0Z_26),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_25),
            .carryout(un1_M_this_warmup_d_cry_26),
            .clk(N__39394),
            .ce(),
            .sr(N__36833));
    defparam M_this_warmup_q_27_LC_10_23_2.C_ON=1'b1;
    defparam M_this_warmup_q_27_LC_10_23_2.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_27_LC_10_23_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 M_this_warmup_q_27_LC_10_23_2 (
            .in0(_gnd_net_),
            .in1(N__16547),
            .in2(_gnd_net_),
            .in3(N__16541),
            .lcout(M_this_warmup_qZ0Z_27),
            .ltout(),
            .carryin(un1_M_this_warmup_d_cry_26),
            .carryout(un1_M_this_warmup_d_cry_27),
            .clk(N__39394),
            .ce(),
            .sr(N__36833));
    defparam M_this_warmup_q_28_LC_10_23_3.C_ON=1'b0;
    defparam M_this_warmup_q_28_LC_10_23_3.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_28_LC_10_23_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 M_this_warmup_q_28_LC_10_23_3 (
            .in0(_gnd_net_),
            .in1(N__16534),
            .in2(_gnd_net_),
            .in3(N__16538),
            .lcout(M_this_warmup_qZ0Z_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39394),
            .ce(),
            .sr(N__36833));
    defparam M_this_status_flags_q_0_LC_10_23_4.C_ON=1'b0;
    defparam M_this_status_flags_q_0_LC_10_23_4.SEQ_MODE=4'b1000;
    defparam M_this_status_flags_q_0_LC_10_23_4.LUT_INIT=16'b1111111110101010;
    LogicCell40 M_this_status_flags_q_0_LC_10_23_4 (
            .in0(N__16535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18831),
            .lcout(M_this_status_flags_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39394),
            .ce(),
            .sr(N__36833));
    defparam M_this_data_tmp_q_esr_8_LC_10_27_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_8_LC_10_27_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_8_LC_10_27_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_8_LC_10_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38103),
            .lcout(M_this_data_tmp_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39411),
            .ce(N__19426),
            .sr(N__36837));
    defparam M_this_data_tmp_q_esr_14_LC_10_27_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_14_LC_10_27_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_14_LC_10_27_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_14_LC_10_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37388),
            .lcout(M_this_data_tmp_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39411),
            .ce(N__19426),
            .sr(N__36837));
    defparam M_this_data_tmp_q_esr_10_LC_10_27_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_10_LC_10_27_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_10_LC_10_27_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_10_LC_10_27_7 (
            .in0(N__37649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39411),
            .ce(N__19426),
            .sr(N__36837));
    defparam \this_start_data_delay.M_last_q_RNILN151_LC_10_28_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNILN151_LC_10_28_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNILN151_LC_10_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNILN151_LC_10_28_0  (
            .in0(_gnd_net_),
            .in1(N__16655),
            .in2(_gnd_net_),
            .in3(N__19328),
            .lcout(M_this_oam_ram_write_data_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINP151_LC_10_28_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINP151_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINP151_LC_10_28_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNINP151_LC_10_28_4  (
            .in0(_gnd_net_),
            .in1(N__17168),
            .in2(_gnd_net_),
            .in3(N__19327),
            .lcout(M_this_oam_ram_write_data_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_7_LC_10_29_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_7_LC_10_29_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_7_LC_10_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_7_LC_10_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38729),
            .lcout(M_this_data_tmp_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39421),
            .ce(N__23621),
            .sr(N__36842));
    defparam M_this_data_tmp_q_esr_5_LC_10_29_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_5_LC_10_29_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_5_LC_10_29_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_5_LC_10_29_7 (
            .in0(N__38918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39421),
            .ce(N__23621),
            .sr(N__36842));
    defparam M_this_data_tmp_q_esr_22_LC_10_30_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_22_LC_10_30_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_22_LC_10_30_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_22_LC_10_30_1 (
            .in0(N__37396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39427),
            .ce(N__21851),
            .sr(N__36845));
    defparam M_this_data_tmp_q_esr_16_LC_10_30_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_16_LC_10_30_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_16_LC_10_30_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_16_LC_10_30_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38101),
            .lcout(M_this_data_tmp_qZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39427),
            .ce(N__21851),
            .sr(N__36845));
    defparam \this_start_data_delay.M_last_q_RNI87IG1_LC_10_31_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI87IG1_LC_10_31_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI87IG1_LC_10_31_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI87IG1_LC_10_31_4  (
            .in0(N__38730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19364),
            .lcout(M_this_oam_ram_write_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINQ251_LC_10_31_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINQ251_LC_10_31_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINQ251_LC_10_31_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNINQ251_LC_10_31_6  (
            .in0(N__19363),
            .in1(N__19844),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_write_data_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIPS251_LC_10_31_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIPS251_LC_10_31_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIPS251_LC_10_31_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIPS251_LC_10_31_7  (
            .in0(_gnd_net_),
            .in1(N__19362),
            .in2(_gnd_net_),
            .in3(N__17774),
            .lcout(M_this_oam_ram_write_data_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_11_7_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_wclke_3_LC_11_7_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_wclke_3_LC_11_7_2  (
            .in0(N__32222),
            .in1(N__32126),
            .in2(N__32036),
            .in3(N__31919),
            .lcout(\this_spr_ram.mem_WE_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_11_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_wclke_3_LC_11_9_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_spr_ram.mem_mem_0_0_wclke_3_LC_11_9_6  (
            .in0(N__32218),
            .in1(N__32125),
            .in2(N__32032),
            .in3(N__31914),
            .lcout(\this_spr_ram.mem_WE_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_5_LC_11_13_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_5_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_5_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_5_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16736),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39310),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_11_14_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_7_0_wclke_3_LC_11_14_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_spr_ram.mem_mem_7_0_wclke_3_LC_11_14_0  (
            .in0(N__32213),
            .in1(N__32118),
            .in2(N__32030),
            .in3(N__31898),
            .lcout(\this_spr_ram.mem_WE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_34_i_LC_11_14_1 .C_ON=1'b0;
    defparam \this_vga_signals.N_34_i_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_34_i_LC_11_14_1 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \this_vga_signals.N_34_i_LC_11_14_1  (
            .in0(N__17892),
            .in1(N__22136),
            .in2(N__18752),
            .in3(N__19628),
            .lcout(N_34_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_14_LC_11_14_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_14_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_14_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_14_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16682),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39316),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI3UQE7_4_LC_11_15_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI3UQE7_4_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI3UQE7_4_LC_11_15_0 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \this_ppu.M_state_q_RNI3UQE7_4_LC_11_15_0  (
            .in0(N__21780),
            .in1(N__21579),
            .in2(N__21374),
            .in3(N__21519),
            .lcout(\this_ppu.M_oam_curr_qc_0_1 ),
            .ltout(\this_ppu.M_oam_curr_qc_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_3_LC_11_15_1 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_3_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_3_LC_11_15_1 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \this_ppu.M_oam_curr_q_3_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__18223),
            .in2(N__16817),
            .in3(N__18274),
            .lcout(M_this_ppu_oam_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39324),
            .ce(),
            .sr(N__38963));
    defparam \this_ppu.M_oam_curr_q_4_LC_11_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_4_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_4_LC_11_15_2 .LUT_INIT=16'b0110110000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_4_LC_11_15_2  (
            .in0(N__18275),
            .in1(N__18650),
            .in2(N__18236),
            .in3(N__18889),
            .lcout(M_this_ppu_oam_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39324),
            .ce(),
            .sr(N__38963));
    defparam \this_ppu.M_oam_curr_q_2_LC_11_15_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_2_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_2_LC_11_15_4 .LUT_INIT=16'b0100100011000000;
    LogicCell40 \this_ppu.M_oam_curr_q_2_LC_11_15_4  (
            .in0(N__18388),
            .in1(N__18888),
            .in2(N__18317),
            .in3(N__18445),
            .lcout(M_this_ppu_oam_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39324),
            .ce(),
            .sr(N__38963));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_4_LC_11_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_4_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_a2_4_LC_11_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_a2_4_LC_11_15_6  (
            .in0(N__18387),
            .in1(N__18304),
            .in2(N__18926),
            .in3(N__18517),
            .lcout(\this_ppu.m35_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_1_LC_11_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_1_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_1_LC_11_16_0 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_1_LC_11_16_0  (
            .in0(N__18392),
            .in1(N__18885),
            .in2(_gnd_net_),
            .in3(N__18444),
            .lcout(M_this_ppu_oam_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39332),
            .ce(),
            .sr(N__38960));
    defparam \this_ppu.M_oam_curr_q_0_LC_11_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_0_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_0_LC_11_16_3 .LUT_INIT=16'b1000001000001010;
    LogicCell40 \this_ppu.M_oam_curr_q_0_LC_11_16_3  (
            .in0(N__18886),
            .in1(N__18570),
            .in2(N__18533),
            .in3(N__18476),
            .lcout(M_this_ppu_oam_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39332),
            .ce(),
            .sr(N__38960));
    defparam \this_ppu.M_screen_x_q_1_LC_11_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_1_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_1_LC_11_17_0 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_screen_x_q_1_LC_11_17_0  (
            .in0(N__17143),
            .in1(N__16965),
            .in2(N__16942),
            .in3(N__16862),
            .lcout(M_this_ppu_vram_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_5_LC_11_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_5_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_5_LC_11_17_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_screen_x_q_5_LC_11_17_1  (
            .in0(N__17016),
            .in1(N__17141),
            .in2(_gnd_net_),
            .in3(N__17036),
            .lcout(M_this_ppu_vram_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_0_LC_11_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_0_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_0_LC_11_17_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_ppu.M_screen_x_q_0_LC_11_17_2  (
            .in0(N__22269),
            .in1(N__30900),
            .in2(N__16941),
            .in3(N__16861),
            .lcout(M_this_ppu_vram_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_11_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIB9B9C_11_LC_11_17_3 .LUT_INIT=16'b0000111011111110;
    LogicCell40 \this_ppu.M_state_q_RNIB9B9C_11_LC_11_17_3  (
            .in0(N__20971),
            .in1(N__21114),
            .in2(N__21166),
            .in3(N__21188),
            .lcout(\this_ppu.N_827_0 ),
            .ltout(\this_ppu.N_827_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_11_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNIM77RC_1_LC_11_17_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNIM77RC_1_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__16964),
            .in2(N__17042),
            .in3(N__16927),
            .lcout(\this_ppu.un1_M_screen_x_q_c2 ),
            .ltout(\this_ppu.un1_M_screen_x_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNIUC1MD_4_LC_11_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNIUC1MD_4_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNIUC1MD_4_LC_11_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNIUC1MD_4_LC_11_17_5  (
            .in0(N__16833),
            .in1(N__16883),
            .in2(N__17039),
            .in3(N__17880),
            .lcout(\this_ppu.un1_M_screen_x_q_c5 ),
            .ltout(\this_ppu.un1_M_screen_x_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_6_LC_11_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_6_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_6_LC_11_17_6 .LUT_INIT=16'b0010100010001000;
    LogicCell40 \this_ppu.M_screen_x_q_6_LC_11_17_6  (
            .in0(N__17142),
            .in1(N__16993),
            .in2(N__17030),
            .in3(N__17017),
            .lcout(M_this_ppu_vram_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_2_LC_11_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_2_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_2_LC_11_17_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \this_ppu.M_screen_x_q_2_LC_11_17_7  (
            .in0(N__30899),
            .in1(N__22270),
            .in2(N__16896),
            .in3(N__16982),
            .lcout(M_this_ppu_vram_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39340),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_RNID854D_1_LC_11_18_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_RNID854D_1_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_x_q_RNID854D_1_LC_11_18_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_screen_x_q_RNID854D_1_LC_11_18_0  (
            .in0(N__16966),
            .in1(N__16928),
            .in2(N__16900),
            .in3(N__16860),
            .lcout(\this_ppu.un1_M_screen_x_q_c3 ),
            .ltout(\this_ppu.un1_M_screen_x_q_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_4_LC_11_18_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_4_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_4_LC_11_18_1 .LUT_INIT=16'b0110110000000000;
    LogicCell40 \this_ppu.M_screen_x_q_4_LC_11_18_1  (
            .in0(N__17885),
            .in1(N__16834),
            .in2(N__16847),
            .in3(N__17144),
            .lcout(M_this_ppu_vram_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39351),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_6_LC_11_18_2 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_6_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_6_LC_11_18_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_6_LC_11_18_2  (
            .in0(N__19160),
            .in1(N__21440),
            .in2(N__30932),
            .in3(N__19025),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39351),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_18_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_18_4  (
            .in0(N__19001),
            .in1(N__28654),
            .in2(_gnd_net_),
            .in3(N__28596),
            .lcout(\this_vga_signals.i22_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_11_18_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIGL6V4_0_LC_11_18_6 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \this_ppu.M_state_q_RNIGL6V4_0_LC_11_18_6  (
            .in0(N__30894),
            .in1(N__21569),
            .in2(_gnd_net_),
            .in3(N__21506),
            .lcout(\this_ppu.N_1210_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_x_q_3_LC_11_18_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_x_q_3_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_x_q_3_LC_11_18_7 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \this_ppu.M_screen_x_q_3_LC_11_18_7  (
            .in0(N__17884),
            .in1(N__30895),
            .in2(N__22274),
            .in3(N__17126),
            .lcout(M_this_ppu_vram_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39351),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_0_LC_11_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_0_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_0_LC_11_19_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_0_LC_11_19_0  (
            .in0(N__21439),
            .in1(N__21209),
            .in2(N__31019),
            .in3(N__19159),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39359),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_13_LC_11_19_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_13_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_13_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_13_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17120),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39359),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_12_LC_11_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_12_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17111),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39359),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_LC_11_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m13_0_a2_LC_11_19_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m13_0_a2_LC_11_19_4  (
            .in0(N__21647),
            .in1(N__21570),
            .in2(_gnd_net_),
            .in3(N__21504),
            .lcout(),
            .ltout(\this_ppu.N_844_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_0_LC_11_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_0_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_0_LC_11_19_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \this_ppu.M_state_q_0_LC_11_19_5  (
            .in0(N__21373),
            .in1(N__17102),
            .in2(N__17093),
            .in3(N__31011),
            .lcout(\this_ppu.M_state_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39359),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_11_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIRJK11_1_LC_11_19_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNIRJK11_1_LC_11_19_7  (
            .in0(N__21113),
            .in1(N__23951),
            .in2(N__20977),
            .in3(N__17083),
            .lcout(\this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_warmup_q_1_LC_11_20_0.C_ON=1'b0;
    defparam M_this_warmup_q_1_LC_11_20_0.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_1_LC_11_20_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 M_this_warmup_q_1_LC_11_20_0 (
            .in0(N__17059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17072),
            .lcout(M_this_warmup_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39368),
            .ce(),
            .sr(N__36828));
    defparam M_this_warmup_q_0_LC_11_20_1.C_ON=1'b0;
    defparam M_this_warmup_q_0_LC_11_20_1.SEQ_MODE=4'b1000;
    defparam M_this_warmup_q_0_LC_11_20_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 M_this_warmup_q_0_LC_11_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17058),
            .lcout(M_this_warmup_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39368),
            .ce(),
            .sr(N__36828));
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_11_20_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIUU07_9_LC_11_20_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIUU07_9_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17528),
            .lcout(\this_ppu.M_oam_cache_read_data_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_11_21_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_11_21_3 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_11_21_3  (
            .in0(N__32670),
            .in1(N__17522),
            .in2(_gnd_net_),
            .in3(N__22737),
            .lcout(M_this_ppu_spr_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI41OT_2_LC_11_22_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI41OT_2_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI41OT_2_LC_11_22_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNI41OT_2_LC_11_22_5  (
            .in0(N__21714),
            .in1(N__20978),
            .in2(N__17270),
            .in3(N__23955),
            .lcout(this_ppu_N_247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_6_LC_11_26_4.C_ON=1'b0;
    defparam M_this_oam_address_q_6_LC_11_26_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_6_LC_11_26_4.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_6_LC_11_26_4 (
            .in0(N__17214),
            .in1(N__25212),
            .in2(_gnd_net_),
            .in3(N__19435),
            .lcout(M_this_oam_address_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39405),
            .ce(),
            .sr(N__38952));
    defparam M_this_oam_address_q_7_LC_11_26_5.C_ON=1'b0;
    defparam M_this_oam_address_q_7_LC_11_26_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_7_LC_11_26_5.LUT_INIT=16'b0000011000001100;
    LogicCell40 M_this_oam_address_q_7_LC_11_26_5 (
            .in0(N__19436),
            .in1(N__17182),
            .in2(N__25217),
            .in3(N__17215),
            .lcout(M_this_oam_address_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39405),
            .ce(),
            .sr(N__38952));
    defparam M_this_data_tmp_q_esr_20_LC_11_27_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_20_LC_11_27_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_20_LC_11_27_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_20_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37466),
            .lcout(M_this_data_tmp_qZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39408),
            .ce(N__21824),
            .sr(N__36835));
    defparam M_this_data_tmp_q_esr_12_LC_11_28_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_12_LC_11_28_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_12_LC_11_28_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_12_LC_11_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37506),
            .lcout(M_this_data_tmp_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39412),
            .ce(N__19427),
            .sr(N__36838));
    defparam M_this_data_tmp_q_esr_15_LC_11_28_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_15_LC_11_28_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_15_LC_11_28_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_15_LC_11_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38768),
            .lcout(M_this_data_tmp_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39412),
            .ce(N__19427),
            .sr(N__36838));
    defparam M_this_data_tmp_q_esr_13_LC_11_28_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_13_LC_11_28_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_13_LC_11_28_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_13_LC_11_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38917),
            .lcout(M_this_data_tmp_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39412),
            .ce(N__19427),
            .sr(N__36838));
    defparam M_this_data_tmp_q_esr_11_LC_11_28_6.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_11_LC_11_28_6.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_11_LC_11_28_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_11_LC_11_28_6 (
            .in0(N__37878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39412),
            .ce(N__19427),
            .sr(N__36838));
    defparam M_this_data_tmp_q_esr_9_LC_11_28_7.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_9_LC_11_28_7.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_9_LC_11_28_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_9_LC_11_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37735),
            .lcout(M_this_data_tmp_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39412),
            .ce(N__19427),
            .sr(N__36838));
    defparam \this_start_data_delay.M_last_q_RNI5KDD1_LC_11_29_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI5KDD1_LC_11_29_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI5KDD1_LC_11_29_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI5KDD1_LC_11_29_1  (
            .in0(N__19298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21869),
            .lcout(M_this_oam_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIMP251_LC_11_29_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIMP251_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIMP251_LC_11_29_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIMP251_LC_11_29_2  (
            .in0(_gnd_net_),
            .in1(N__19297),
            .in2(_gnd_net_),
            .in3(N__17615),
            .lcout(M_this_oam_ram_write_data_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI6LDD1_LC_11_29_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI6LDD1_LC_11_29_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI6LDD1_LC_11_29_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI6LDD1_LC_11_29_3  (
            .in0(N__19299),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19850),
            .lcout(M_this_oam_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIDSDD1_LC_11_29_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIDSDD1_LC_11_29_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIDSDD1_LC_11_29_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIDSDD1_LC_11_29_5  (
            .in0(N__19301),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17582),
            .lcout(M_this_oam_ram_write_data_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI8NDD1_LC_11_29_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI8NDD1_LC_11_29_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI8NDD1_LC_11_29_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI8NDD1_LC_11_29_6  (
            .in0(_gnd_net_),
            .in1(N__19296),
            .in2(_gnd_net_),
            .in3(N__19208),
            .lcout(M_this_oam_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIMO151_LC_11_29_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIMO151_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIMO151_LC_11_29_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIMO151_LC_11_29_7  (
            .in0(N__19300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17555),
            .lcout(M_this_oam_ram_write_data_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_17_LC_11_30_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_17_LC_11_30_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_17_LC_11_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_17_LC_11_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37734),
            .lcout(M_this_data_tmp_qZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39422),
            .ce(N__21850),
            .sr(N__36843));
    defparam M_this_data_tmp_q_esr_23_LC_11_30_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_23_LC_11_30_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_23_LC_11_30_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_23_LC_11_30_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38769),
            .lcout(M_this_data_tmp_qZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39422),
            .ce(N__21850),
            .sr(N__36843));
    defparam \this_start_data_delay.M_last_q_RNIU0251_LC_11_31_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIU0251_LC_11_31_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIU0251_LC_11_31_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIU0251_LC_11_31_2  (
            .in0(_gnd_net_),
            .in1(N__21860),
            .in2(_gnd_net_),
            .in3(N__19384),
            .lcout(M_this_oam_ram_write_data_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI54IG1_LC_11_31_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI54IG1_LC_11_31_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI54IG1_LC_11_31_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI54IG1_LC_11_31_3  (
            .in0(N__19386),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37507),
            .lcout(M_this_oam_ram_write_data_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI21IG1_LC_11_31_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI21IG1_LC_11_31_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI21IG1_LC_11_31_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI21IG1_LC_11_31_6  (
            .in0(_gnd_net_),
            .in1(N__37715),
            .in2(_gnd_net_),
            .in3(N__19385),
            .lcout(M_this_oam_ram_write_data_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_12_9_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_12_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_12_9_4  (
            .in0(N__20825),
            .in1(N__17738),
            .in2(_gnd_net_),
            .in3(N__17723),
            .lcout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_12_10_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_12_10_0 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_12_10_0  (
            .in0(N__19925),
            .in1(N__17936),
            .in2(N__19693),
            .in3(N__17711),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_12_10_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_12_10_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_12_10_1  (
            .in0(N__19926),
            .in1(N__17633),
            .in2(N__17705),
            .in3(N__17672),
            .lcout(M_this_spr_ram_read_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_12_10_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_12_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_12_10_5  (
            .in0(N__17702),
            .in1(N__17684),
            .in2(_gnd_net_),
            .in3(N__20839),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_12_10_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_12_10_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_12_10_6  (
            .in0(N__20840),
            .in1(N__17666),
            .in2(_gnd_net_),
            .in3(N__17651),
            .lcout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_12_11_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_12_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_12_11_2  (
            .in0(N__20826),
            .in1(N__17972),
            .in2(_gnd_net_),
            .in3(N__17954),
            .lcout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_12_11_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_12_11_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_12_11_6  (
            .in0(N__20827),
            .in1(N__17930),
            .in2(_gnd_net_),
            .in3(N__17915),
            .lcout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_12_12_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_12_LC_12_12_3 .LUT_INIT=16'b0001101000011111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_12_LC_12_12_3  (
            .in0(N__19906),
            .in1(N__19967),
            .in2(N__19694),
            .in3(N__17903),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.m21_LC_12_13_1 .C_ON=1'b0;
    defparam \this_vga_signals.m21_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.m21_LC_12_13_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.m21_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__17896),
            .in2(_gnd_net_),
            .in3(N__22135),
            .lcout(\this_vga_signals.N_22_0 ),
            .ltout(\this_vga_signals.N_22_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_856_i_LC_12_13_2 .C_ON=1'b0;
    defparam \this_vga_signals.N_856_i_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_856_i_LC_12_13_2 .LUT_INIT=16'b1010111000000100;
    LogicCell40 \this_vga_signals.N_856_i_LC_12_13_2  (
            .in0(N__18748),
            .in1(N__22075),
            .in2(N__17849),
            .in3(N__18611),
            .lcout(N_856_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_12_13_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_12_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_12_13_3  (
            .in0(N__17831),
            .in1(N__17813),
            .in2(_gnd_net_),
            .in3(N__20863),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_12_13_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_11_LC_12_13_4 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_11_LC_12_13_4  (
            .in0(N__20780),
            .in1(N__19910),
            .in2(N__17798),
            .in3(N__17795),
            .lcout(M_this_spr_ram_read_data_3),
            .ltout(M_this_spr_ram_read_data_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_25_0_i_LC_12_13_5 .C_ON=1'b0;
    defparam \this_vga_signals.N_25_0_i_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_25_0_i_LC_12_13_5 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \this_vga_signals.N_25_0_i_LC_12_13_5  (
            .in0(N__18747),
            .in1(N__18706),
            .in2(N__17789),
            .in3(N__22361),
            .lcout(N_25_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_12_13_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_12_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18161),
            .lcout(\this_ppu.M_oam_cache_read_data_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_12_14_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_12_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_12_14_3  (
            .in0(N__20852),
            .in1(N__18155),
            .in2(_gnd_net_),
            .in3(N__18137),
            .lcout(\this_spr_ram.mem_mem_0_1_RNIM6VFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_12_14_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII6H51_6_LC_12_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_RNII6H51_6_LC_12_14_5  (
            .in0(N__21163),
            .in1(N__20767),
            .in2(N__21778),
            .in3(N__22042),
            .lcout(\this_ppu.M_state_q_inv_1 ),
            .ltout(\this_ppu.M_state_q_inv_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_12_LC_12_14_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_12_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_12_LC_12_14_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \this_spr_ram.mem_radreg_12_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__18125),
            .in2(N__18113),
            .in3(N__18110),
            .lcout(\this_spr_ram.mem_radregZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39311),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_5_LC_12_15_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_5_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_5_LC_12_15_0 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \this_ppu.M_state_q_5_LC_12_15_0  (
            .in0(N__18571),
            .in1(N__21376),
            .in2(N__18089),
            .in3(N__30983),
            .lcout(\this_ppu.M_state_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39317),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_12_15_1 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_12_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_12_15_1  (
            .in0(N__18077),
            .in1(N__18059),
            .in2(_gnd_net_),
            .in3(N__20865),
            .lcout(\this_spr_ram.mem_mem_1_1_RNIOA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_12_15_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_LC_12_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_LC_12_15_2  (
            .in0(N__20866),
            .in1(N__18044),
            .in2(_gnd_net_),
            .in3(N__18029),
            .lcout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_12_15_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_12_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_12_15_3  (
            .in0(N__18011),
            .in1(N__20864),
            .in2(_gnd_net_),
            .in3(N__17993),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_12_15_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_12_15_4 .LUT_INIT=16'b0010011000110111;
    LogicCell40 \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_12_15_4  (
            .in0(N__19915),
            .in1(N__19682),
            .in2(N__17981),
            .in3(N__17978),
            .lcout(),
            .ltout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_12_15_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_12_15_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_12_15_5  (
            .in0(N__19927),
            .in1(N__18767),
            .in2(N__18761),
            .in3(N__18758),
            .lcout(M_this_spr_ram_read_data_2),
            .ltout(M_this_spr_ram_read_data_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.N_28_0_i_LC_12_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.N_28_0_i_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.N_28_0_i_LC_12_15_6 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \this_vga_signals.N_28_0_i_LC_12_15_6  (
            .in0(N__18746),
            .in1(N__18710),
            .in2(N__18695),
            .in3(N__22397),
            .lcout(N_28_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIGIC2L_4_LC_12_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIGIC2L_4_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIGIC2L_4_LC_12_16_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIGIC2L_4_LC_12_16_0  (
            .in0(N__18646),
            .in1(N__18221),
            .in2(_gnd_net_),
            .in3(N__18273),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_d25_LC_12_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_d25_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_d25_LC_12_16_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_oam_curr_d25_LC_12_16_1  (
            .in0(N__18617),
            .in1(N__18610),
            .in2(N__18596),
            .in3(N__19627),
            .lcout(\this_ppu.M_oam_curr_dZ0Z25 ),
            .ltout(\this_ppu.M_oam_curr_dZ0Z25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIQ09CG_6_LC_12_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIQ09CG_6_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIQ09CG_6_LC_12_16_2 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \this_ppu.M_state_q_RNIQ09CG_6_LC_12_16_2  (
            .in0(N__22041),
            .in1(N__21165),
            .in2(N__18581),
            .in3(N__22015),
            .lcout(\this_ppu.N_834_0 ),
            .ltout(\this_ppu.N_834_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNIEH7HK_0_LC_12_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNIEH7HK_0_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNIEH7HK_0_LC_12_16_3 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \this_ppu.M_oam_curr_q_RNIEH7HK_0_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__18513),
            .in2(N__18479),
            .in3(N__18475),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c1 ),
            .ltout(\this_ppu.un1_M_oam_curr_q_1_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNITVPPK_2_LC_12_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNITVPPK_2_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNITVPPK_2_LC_12_16_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNITVPPK_2_LC_12_16_4  (
            .in0(N__18386),
            .in1(_gnd_net_),
            .in2(N__18353),
            .in3(N__18303),
            .lcout(\this_ppu.un1_M_oam_curr_q_1_c3 ),
            .ltout(\this_ppu.un1_M_oam_curr_q_1_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_RNI5CAKS_3_LC_12_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_RNI5CAKS_3_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_oam_curr_q_RNI5CAKS_3_LC_12_16_5 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_RNI5CAKS_3_LC_12_16_5  (
            .in0(N__18222),
            .in1(_gnd_net_),
            .in2(N__18188),
            .in3(N__18787),
            .lcout(\this_ppu.N_778_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_oam_curr_q_5_LC_12_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_5_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_5_LC_12_16_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \this_ppu.M_oam_curr_q_5_LC_12_16_6  (
            .in0(N__18927),
            .in1(N__18887),
            .in2(_gnd_net_),
            .in3(N__18955),
            .lcout(M_this_ppu_oam_addr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39325),
            .ce(),
            .sr(N__38957));
    defparam \this_ppu.M_oam_curr_q_6_LC_12_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_oam_curr_q_6_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_oam_curr_q_6_LC_12_16_7 .LUT_INIT=16'b0110110000000000;
    LogicCell40 \this_ppu.M_oam_curr_q_6_LC_12_16_7  (
            .in0(N__18956),
            .in1(N__18859),
            .in2(N__18928),
            .in3(N__18890),
            .lcout(\this_ppu.M_oam_curr_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39325),
            .ce(),
            .sr(N__38957));
    defparam \this_ppu.M_state_q_7_LC_12_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_7_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_7_LC_12_17_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_ppu.M_state_q_7_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__30990),
            .in2(_gnd_net_),
            .in3(N__22019),
            .lcout(\this_ppu.M_state_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_10_LC_12_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_10_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_10_LC_12_17_1 .LUT_INIT=16'b0000111100000010;
    LogicCell40 \this_ppu.M_state_q_10_LC_12_17_1  (
            .in0(N__22250),
            .in1(N__18845),
            .in2(N__36963),
            .in3(N__20976),
            .lcout(\this_ppu.M_state_qZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_15_LC_12_17_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_15_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_15_LC_12_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_15_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18812),
            .lcout(\this_ppu.M_oam_cache_read_data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39333),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIF37M7_4_LC_12_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIF37M7_4_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIF37M7_4_LC_12_17_6 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \this_ppu.M_state_q_RNIF37M7_4_LC_12_17_6  (
            .in0(N__21779),
            .in1(N__36929),
            .in2(N__21359),
            .in3(N__22249),
            .lcout(\this_ppu.N_784_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_12_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNO_0_1_LC_12_18_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNO_0_1_LC_12_18_0  (
            .in0(N__18979),
            .in1(N__28655),
            .in2(_gnd_net_),
            .in3(N__28612),
            .lcout(),
            .ltout(\this_vga_signals.N_859_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_1_LC_12_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_1_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_1_LC_12_18_1 .LUT_INIT=16'b0111010011001100;
    LogicCell40 \this_vga_signals.M_lcounter_q_1_LC_12_18_1  (
            .in0(N__28614),
            .in1(N__19000),
            .in2(N__18776),
            .in3(N__29778),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_12_18_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI94M7_13_LC_12_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI94M7_13_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18773),
            .lcout(\this_ppu.M_oam_cache_read_data_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_5_LC_12_18_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_5_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_5_LC_12_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m9_0_a2_5_LC_12_18_3  (
            .in0(N__19090),
            .in1(N__19066),
            .in2(N__19042),
            .in3(N__19114),
            .lcout(),
            .ltout(\this_ppu.m9_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_LC_12_18_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_LC_12_18_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m9_0_a2_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19010),
            .in3(N__21242),
            .lcout(\this_ppu.N_97_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_0_LC_12_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_0_LC_12_18_6 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_lcounter_q_0_LC_12_18_6 .LUT_INIT=16'b0100101011101010;
    LogicCell40 \this_vga_signals.M_lcounter_q_0_LC_12_18_6  (
            .in0(N__18980),
            .in1(N__19007),
            .in2(N__29791),
            .in3(N__28613),
            .lcout(\this_vga_signals.M_lcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39341),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_12_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_12_18_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_12_18_7  (
            .in0(N__18996),
            .in1(N__18978),
            .in2(_gnd_net_),
            .in3(N__35276),
            .lcout(N_52_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNI58DK1_5_LC_12_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNI58DK1_5_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNI58DK1_5_LC_12_19_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_ppu.M_state_q_RNI58DK1_5_LC_12_19_0  (
            .in0(N__21164),
            .in1(N__20771),
            .in2(_gnd_net_),
            .in3(N__18968),
            .lcout(\this_ppu.N_814 ),
            .ltout(\this_ppu.N_814_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIOVN89_10_LC_12_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIOVN89_10_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIOVN89_10_LC_12_19_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_state_q_RNIOVN89_10_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(N__21341),
            .in2(N__18962),
            .in3(N__21949),
            .lcout(\this_ppu.N_806 ),
            .ltout(\this_ppu.N_806_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_2_LC_12_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_2_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_2_LC_12_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_2_LC_12_19_2  (
            .in0(N__30995),
            .in1(N__21435),
            .in2(N__18959),
            .in3(N__19124),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_5_LC_12_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_5_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_5_LC_12_19_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_5_LC_12_19_3  (
            .in0(N__21438),
            .in1(N__19158),
            .in2(N__31018),
            .in3(N__19055),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_3_LC_12_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_3_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_3_LC_12_19_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_3_LC_12_19_4  (
            .in0(N__19156),
            .in1(N__21436),
            .in2(N__31015),
            .in3(N__19103),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_4_LC_12_19_6 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_4_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_4_LC_12_19_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_4_LC_12_19_6  (
            .in0(N__19157),
            .in1(N__21437),
            .in2(N__31016),
            .in3(N__19079),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_1_LC_12_19_7 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_1_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_1_LC_12_19_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_1_LC_12_19_7  (
            .in0(N__21434),
            .in1(N__19155),
            .in2(N__31017),
            .in3(N__19133),
            .lcout(\this_ppu.M_pixel_cnt_qZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39352),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_LC_12_20_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_LC_12_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__21668),
            .in2(N__21235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_1_LC_12_20_1 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_1_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_1_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__21791),
            .in2(N__21278),
            .in3(N__19127),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_0 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_2_LC_12_20_2 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_2_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_2_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_2_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__21803),
            .in2(N__21296),
            .in3(N__19118),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_1 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_3_LC_12_20_3 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_3_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_3_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_3_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__19115),
            .in2(N__21908),
            .in3(N__19097),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_2 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_4_LC_12_20_4 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_4_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_4_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_4_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__19199),
            .in2(N__19094),
            .in3(N__19073),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_3 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_5_LC_12_20_5 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_5_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_5_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_5_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__19166),
            .in2(N__19070),
            .in3(N__19049),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_4 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_6_LC_12_20_6 .C_ON=1'b1;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_6_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_6_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__21797),
            .in2(N__19046),
            .in3(N__19013),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_pixel_cnt_q_1_cry_5 ),
            .carryout(\this_ppu.un1_M_pixel_cnt_q_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_12_20_7 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_12_20_7 .LUT_INIT=16'b1000011101111000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_12_20_7  (
            .in0(N__21991),
            .in1(N__21950),
            .in2(N__21262),
            .in3(N__19202),
            .lcout(\this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_1_10_LC_12_21_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_1_10_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_1_10_LC_12_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_1_10_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__21994),
            .in2(_gnd_net_),
            .in3(N__21947),
            .lcout(\this_ppu.M_state_q_RNISP3R6_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_21_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__19193),
            .in2(_gnd_net_),
            .in3(N__23995),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_10_LC_12_21_7 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_10_LC_12_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_10_LC_12_21_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_10_LC_12_21_7  (
            .in0(N__21948),
            .in1(_gnd_net_),
            .in2(N__21998),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_state_q_RNISP3R6Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_0_LC_12_24_4.C_ON=1'b0;
    defparam M_this_oam_address_q_0_LC_12_24_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_0_LC_12_24_4.LUT_INIT=16'b0000010100001010;
    LogicCell40 M_this_oam_address_q_0_LC_12_24_4 (
            .in0(N__23658),
            .in1(_gnd_net_),
            .in2(N__25198),
            .in3(N__23704),
            .lcout(M_this_oam_address_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39391),
            .ce(),
            .sr(N__38954));
    defparam M_this_oam_address_q_3_LC_12_25_0.C_ON=1'b0;
    defparam M_this_oam_address_q_3_LC_12_25_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_3_LC_12_25_0.LUT_INIT=16'b0000000001111000;
    LogicCell40 M_this_oam_address_q_3_LC_12_25_0 (
            .in0(N__21898),
            .in1(N__19552),
            .in2(N__19594),
            .in3(N__25209),
            .lcout(M_this_oam_address_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39395),
            .ce(),
            .sr(N__38953));
    defparam M_this_oam_address_q_4_LC_12_25_3.C_ON=1'b0;
    defparam M_this_oam_address_q_4_LC_12_25_3.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_4_LC_12_25_3.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_4_LC_12_25_3 (
            .in0(N__19461),
            .in1(N__25200),
            .in2(_gnd_net_),
            .in3(N__19528),
            .lcout(M_this_oam_address_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39395),
            .ce(),
            .sr(N__38953));
    defparam M_this_oam_address_q_5_LC_12_25_4.C_ON=1'b0;
    defparam M_this_oam_address_q_5_LC_12_25_4.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_5_LC_12_25_4.LUT_INIT=16'b0000000001101100;
    LogicCell40 M_this_oam_address_q_5_LC_12_25_4 (
            .in0(N__19529),
            .in1(N__19504),
            .in2(N__19468),
            .in3(N__25210),
            .lcout(M_this_oam_address_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39395),
            .ce(),
            .sr(N__38953));
    defparam M_this_oam_address_q_2_LC_12_25_5.C_ON=1'b0;
    defparam M_this_oam_address_q_2_LC_12_25_5.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_2_LC_12_25_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_oam_address_q_2_LC_12_25_5 (
            .in0(N__19551),
            .in1(N__25199),
            .in2(_gnd_net_),
            .in3(N__21897),
            .lcout(M_this_oam_address_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39395),
            .ce(),
            .sr(N__38953));
    defparam M_this_oam_address_q_RNILNG41_3_LC_12_26_1.C_ON=1'b0;
    defparam M_this_oam_address_q_RNILNG41_3_LC_12_26_1.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNILNG41_3_LC_12_26_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 M_this_oam_address_q_RNILNG41_3_LC_12_26_1 (
            .in0(N__21899),
            .in1(N__19587),
            .in2(_gnd_net_),
            .in3(N__19550),
            .lcout(un1_M_this_oam_address_q_c4),
            .ltout(un1_M_this_oam_address_q_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIOKR51_5_LC_12_26_2.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_12_26_2.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIOKR51_5_LC_12_26_2.LUT_INIT=16'b1100000000000000;
    LogicCell40 M_this_oam_address_q_RNIOKR51_5_LC_12_26_2 (
            .in0(_gnd_net_),
            .in1(N__19503),
            .in2(N__19484),
            .in3(N__19460),
            .lcout(un1_M_this_oam_address_q_c6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_12_27_7.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_12_27_7.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_0_1_LC_12_27_7.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_0_1_LC_12_27_7 (
            .in0(N__23758),
            .in1(N__23721),
            .in2(N__23671),
            .in3(N__36947),
            .lcout(N_1240_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIMU531_LC_12_28_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIMU531_LC_12_28_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIMU531_LC_12_28_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIMU531_LC_12_28_0  (
            .in0(N__23763),
            .in1(N__23662),
            .in2(_gnd_net_),
            .in3(N__23719),
            .lcout(M_this_oam_ram_write_data_0_sqmuxa),
            .ltout(M_this_oam_ram_write_data_0_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI32IG1_LC_12_28_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI32IG1_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI32IG1_LC_12_28_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI32IG1_LC_12_28_1  (
            .in0(N__37650),
            .in1(_gnd_net_),
            .in2(N__19409),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_write_data_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_LC_12_28_2.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_12_28_2.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_LC_12_28_2.LUT_INIT=16'b1111001011110000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_LC_12_28_2 (
            .in0(N__23764),
            .in1(N__23720),
            .in2(N__36965),
            .in3(N__23663),
            .lcout(N_1232_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI4JDD1_LC_12_28_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI4JDD1_LC_12_28_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI4JDD1_LC_12_28_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI4JDD1_LC_12_28_3  (
            .in0(N__19214),
            .in1(N__19266),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_oam_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_tmp_q_esr_0_LC_12_29_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_0_LC_12_29_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_0_LC_12_29_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_0_LC_12_29_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38078),
            .lcout(M_this_data_tmp_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39413),
            .ce(N__23619),
            .sr(N__36839));
    defparam M_this_data_tmp_q_esr_4_LC_12_29_1.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_4_LC_12_29_1.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_4_LC_12_29_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_4_LC_12_29_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37522),
            .lcout(M_this_data_tmp_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39413),
            .ce(N__23619),
            .sr(N__36839));
    defparam M_this_data_tmp_q_esr_2_LC_12_29_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_2_LC_12_29_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_2_LC_12_29_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_2_LC_12_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37615),
            .lcout(M_this_data_tmp_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39413),
            .ce(N__23619),
            .sr(N__36839));
    defparam M_this_data_tmp_q_esr_21_LC_12_31_0.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_21_LC_12_31_0.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_21_LC_12_31_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_21_LC_12_31_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38894),
            .lcout(M_this_data_tmp_qZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39423),
            .ce(N__21848),
            .sr(N__36844));
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_13_9_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_13_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_13_9_0  (
            .in0(N__19835),
            .in1(N__19811),
            .in2(_gnd_net_),
            .in3(N__20830),
            .lcout(\this_spr_ram.mem_mem_3_0_RNIQI5GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_9_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_9_2  (
            .in0(N__20824),
            .in1(N__19793),
            .in2(_gnd_net_),
            .in3(N__19778),
            .lcout(\this_spr_ram.mem_mem_0_0_RNIK6VFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_13_9_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_13_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_13_9_4  (
            .in0(N__19763),
            .in1(N__19742),
            .in2(_gnd_net_),
            .in3(N__20829),
            .lcout(\this_spr_ram.mem_mem_1_0_RNIMA1GZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_13_9_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_13_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_13_9_5  (
            .in0(N__20828),
            .in1(N__19727),
            .in2(_gnd_net_),
            .in3(N__19709),
            .lcout(),
            .ltout(\this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_13_9_6 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_13_9_6 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_13_9_6  (
            .in0(N__19692),
            .in1(N__19911),
            .in2(N__19655),
            .in3(N__19652),
            .lcout(\this_spr_ram.mem_DOUT_7_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_13_10_2 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_13_10_2 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_13_10_2  (
            .in0(N__19646),
            .in1(N__19640),
            .in2(N__19928),
            .in3(N__19634),
            .lcout(M_this_spr_ram_read_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_13_LC_13_10_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_13_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_13_LC_13_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_radreg_13_LC_13_10_5  (
            .in0(N__20705),
            .in1(N__20690),
            .in2(_gnd_net_),
            .in3(N__32688),
            .lcout(\this_spr_ram.mem_radregZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39289),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_11_0 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_11_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_11_0  (
            .in0(N__20681),
            .in1(N__20669),
            .in2(_gnd_net_),
            .in3(N__32664),
            .lcout(M_this_ppu_spr_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_11_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_11_2  (
            .in0(N__20441),
            .in1(N__20429),
            .in2(_gnd_net_),
            .in3(N__32663),
            .lcout(M_this_ppu_spr_addr_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_13_11_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_13_11_4 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_13_11_4  (
            .in0(N__32665),
            .in1(N__24927),
            .in2(N__26567),
            .in3(N__24928),
            .lcout(M_this_ppu_spr_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_13_11_7 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_13_11_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_13_11_7  (
            .in0(N__20838),
            .in1(N__19997),
            .in2(_gnd_net_),
            .in3(N__19982),
            .lcout(\this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_radreg_11_LC_13_12_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_radreg_11_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \this_spr_ram.mem_radreg_11_LC_13_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_spr_ram.mem_radreg_11_LC_13_12_5  (
            .in0(N__19961),
            .in1(N__19949),
            .in2(_gnd_net_),
            .in3(N__32669),
            .lcout(\this_spr_ram.mem_radregZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39297),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_4_LC_13_13_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_4_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_4_LC_13_13_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_4_LC_13_13_0  (
            .in0(N__23182),
            .in1(N__22076),
            .in2(_gnd_net_),
            .in3(N__22151),
            .lcout(this_ppu_M_screen_y_q_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39301),
            .ce(N__23060),
            .sr(N__36826));
    defparam \this_ppu.M_state_q_8_LC_13_14_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_8_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_8_LC_13_14_5 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \this_ppu.M_state_q_8_LC_13_14_5  (
            .in0(N__19856),
            .in1(N__36958),
            .in2(N__20741),
            .in3(N__20770),
            .lcout(\this_ppu.M_state_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39306),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_m2_LC_13_15_0 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_m2_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m71_i_m2_LC_13_15_0 .LUT_INIT=16'b1100110011111011;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m71_i_m2_LC_13_15_0  (
            .in0(N__21375),
            .in1(N__21772),
            .in2(N__24049),
            .in3(N__20768),
            .lcout(\this_ppu.N_797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIFCA89_2_LC_13_15_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIFCA89_2_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIFCA89_2_LC_13_15_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIFCA89_2_LC_13_15_1  (
            .in0(N__23096),
            .in1(N__22119),
            .in2(_gnd_net_),
            .in3(N__22096),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c4 ),
            .ltout(\this_ppu.un3_M_screen_y_d_0_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIMH2E9_5_LC_13_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIMH2E9_5_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIMH2E9_5_LC_13_15_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIMH2E9_5_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__22385),
            .in2(N__20915),
            .in3(N__22085),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_4_LC_13_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_4_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_4_LC_13_15_3 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \this_ppu.M_state_q_4_LC_13_15_3  (
            .in0(N__30984),
            .in1(N__21099),
            .in2(N__20912),
            .in3(N__20996),
            .lcout(\this_ppu.M_state_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39312),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_13_15_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_13_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_13_15_4  (
            .in0(N__20897),
            .in1(N__20882),
            .in2(_gnd_net_),
            .in3(N__20867),
            .lcout(\this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_6_LC_13_15_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_6_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_6_LC_13_15_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_state_q_6_LC_13_15_5  (
            .in0(N__20769),
            .in1(N__20737),
            .in2(_gnd_net_),
            .in3(N__36956),
            .lcout(\this_ppu.M_state_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39312),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_9_LC_13_15_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_9_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_state_q_9_LC_13_15_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_ppu.M_state_q_9_LC_13_15_6  (
            .in0(N__36955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20714),
            .lcout(\this_ppu.M_state_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39312),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_13_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_6_LC_13_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_6_LC_13_16_0  (
            .in0(N__24244),
            .in1(N__24164),
            .in2(N__21020),
            .in3(N__24305),
            .lcout(),
            .ltout(\this_ppu.un1_M_surface_x_q_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_6_LC_13_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_6_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_6_LC_13_16_1 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \this_ppu.M_surface_x_q_6_LC_13_16_1  (
            .in0(N__24086),
            .in1(N__22266),
            .in2(N__20708),
            .in3(N__21035),
            .lcout(M_this_ppu_map_addr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39318),
            .ce(),
            .sr(N__36819));
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_o2_LC_13_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_o2_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m35_i_o2_LC_13_16_2 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m35_i_o2_LC_13_16_2  (
            .in0(N__21170),
            .in1(N__21189),
            .in2(_gnd_net_),
            .in3(N__21091),
            .lcout(\this_ppu.N_798_0 ),
            .ltout(\this_ppu.N_798_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_13_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_13_16_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_13_16_3  (
            .in0(N__24574),
            .in1(N__24864),
            .in2(N__21023),
            .in3(N__24914),
            .lcout(\this_ppu.un1_M_surface_x_q_c3 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_3_LC_13_16_4 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_3_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_3_LC_13_16_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \this_ppu.M_surface_x_q_3_LC_13_16_4  (
            .in0(N__21050),
            .in1(N__22267),
            .in2(N__21011),
            .in3(N__24306),
            .lcout(M_this_ppu_map_addr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39318),
            .ce(),
            .sr(N__36819));
    defparam \this_ppu.M_surface_x_q_0_LC_13_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_0_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_0_LC_13_16_6 .LUT_INIT=16'b1111000010011001;
    LogicCell40 \this_ppu.M_surface_x_q_0_LC_13_16_6  (
            .in0(N__24915),
            .in1(N__21008),
            .in2(N__21398),
            .in3(N__22268),
            .lcout(\this_ppu.offset_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39318),
            .ce(),
            .sr(N__36819));
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_13_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_7_LC_13_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_7_LC_13_16_7  (
            .in0(N__22285),
            .in1(N__24163),
            .in2(N__24093),
            .in3(N__24243),
            .lcout(\this_ppu.un1_M_surface_x_q_ac0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_13_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNINHSUC_1_LC_13_17_0 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNINHSUC_1_LC_13_17_0  (
            .in0(N__24863),
            .in1(N__20992),
            .in2(N__21116),
            .in3(N__24913),
            .lcout(\this_ppu.un1_M_surface_x_q_c2 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_13_17_1 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNO_0_5_LC_13_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNO_0_5_LC_13_17_1  (
            .in0(N__24304),
            .in1(N__24245),
            .in2(N__21002),
            .in3(N__24572),
            .lcout(),
            .ltout(\this_ppu.un1_M_surface_x_q_c5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_5_LC_13_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_5_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_5_LC_13_17_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \this_ppu.M_surface_x_q_5_LC_13_17_2  (
            .in0(N__21041),
            .in1(N__22252),
            .in2(N__20999),
            .in3(N__24165),
            .lcout(M_this_ppu_map_addr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39326),
            .ce(),
            .sr(N__36816));
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_13_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNII1FQB_7_LC_13_17_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_ppu.M_state_q_RNII1FQB_7_LC_13_17_3  (
            .in0(N__21155),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21190),
            .lcout(\this_ppu.N_800 ),
            .ltout(\this_ppu.N_800_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_13_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNICH7OC_11_LC_13_17_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \this_ppu.M_state_q_RNICH7OC_11_LC_13_17_4  (
            .in0(N__21112),
            .in1(N__26690),
            .in2(N__20981),
            .in3(N__20975),
            .lcout(N_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_2_LC_13_17_5 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_2_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_2_LC_13_17_5 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_surface_x_q_2_LC_13_17_5  (
            .in0(N__22251),
            .in1(N__21197),
            .in2(N__21062),
            .in3(N__24573),
            .lcout(\this_ppu.M_surface_x_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39326),
            .ce(),
            .sr(N__36816));
    defparam \this_ppu.M_state_q_RNIOVBHC_7_LC_13_17_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIOVBHC_7_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIOVBHC_7_LC_13_17_6 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \this_ppu.M_state_q_RNIOVBHC_7_LC_13_17_6  (
            .in0(N__21191),
            .in1(N__21156),
            .in2(N__21115),
            .in3(N__24912),
            .lcout(\this_ppu.un1_M_surface_x_q_c1 ),
            .ltout(\this_ppu.un1_M_surface_x_q_c1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_13_17_7 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_13_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_13_17_7  (
            .in0(N__24303),
            .in1(N__24571),
            .in2(N__21065),
            .in3(N__24862),
            .lcout(\this_ppu.un1_M_surface_x_q_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_10_LC_13_18_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_10_LC_13_18_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_10_LC_13_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_10_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37652),
            .lcout(M_this_scroll_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_11_LC_13_18_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_11_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_11_LC_13_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_11_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37898),
            .lcout(M_this_scroll_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_12_LC_13_18_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_12_LC_13_18_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_12_LC_13_18_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_12_LC_13_18_2 (
            .in0(N__37529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_13_LC_13_18_3.C_ON=1'b0;
    defparam M_this_scroll_q_esr_13_LC_13_18_3.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_13_LC_13_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_13_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38910),
            .lcout(M_this_scroll_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_14_LC_13_18_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_14_LC_13_18_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_14_LC_13_18_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_14_LC_13_18_4 (
            .in0(N__37352),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_15_LC_13_18_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_15_LC_13_18_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_15_LC_13_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_15_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38760),
            .lcout(M_this_scroll_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_8_LC_13_18_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_8_LC_13_18_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_8_LC_13_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_8_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38129),
            .lcout(M_this_scroll_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam M_this_scroll_q_esr_9_LC_13_18_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_9_LC_13_18_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_9_LC_13_18_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_9_LC_13_18_7 (
            .in0(N__37739),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39334),
            .ce(N__23501),
            .sr(N__36820));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFICF2_5_LC_13_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFICF2_5_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIFICF2_5_LC_13_19_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIFICF2_5_LC_13_19_1  (
            .in0(N__33172),
            .in1(N__23531),
            .in2(_gnd_net_),
            .in3(N__33942),
            .lcout(),
            .ltout(N_829_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m14_0_o2_LC_13_19_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m14_0_o2_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m14_0_o2_LC_13_19_2 .LUT_INIT=16'b1100100000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m14_0_o2_LC_13_19_2  (
            .in0(N__34073),
            .in1(N__34650),
            .in2(N__21383),
            .in3(N__34752),
            .lcout(N_58_0),
            .ltout(N_58_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_13_19_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_13_19_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_13_19_3  (
            .in0(N__29810),
            .in1(N__21594),
            .in2(N__21380),
            .in3(N__29847),
            .lcout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0 ),
            .ltout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_7_LC_13_19_4 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_7_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_pixel_cnt_q_7_LC_13_19_4 .LUT_INIT=16'b1011101110110000;
    LogicCell40 \this_ppu.M_pixel_cnt_q_7_LC_13_19_4  (
            .in0(N__21643),
            .in1(N__21372),
            .in2(N__21305),
            .in3(N__21302),
            .lcout(\this_ppu.M_pixel_cnt_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39342),
            .ce(),
            .sr(N__36822));
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_4_LC_13_19_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_4_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m9_0_a2_4_LC_13_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m9_0_a2_4_LC_13_19_5  (
            .in0(N__21295),
            .in1(N__21274),
            .in2(N__21263),
            .in3(N__21231),
            .lcout(\this_ppu.m9_0_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_0_LC_13_20_0 .C_ON=1'b0;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_0_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_pixel_cnt_q_RNO_0_0_LC_13_20_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_pixel_cnt_q_RNO_0_0_LC_13_20_0  (
            .in0(N__21980),
            .in1(N__21236),
            .in2(_gnd_net_),
            .in3(N__21945),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_13_20_1 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNIJ1SE_10_LC_13_20_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_ppu.M_state_q_RNIJ1SE_10_LC_13_20_1  (
            .in0(N__21710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21777),
            .lcout(\this_ppu.N_60_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_2_10_LC_13_20_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_2_10_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_2_10_LC_13_20_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_2_10_LC_13_20_2  (
            .in0(N__21978),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21943),
            .lcout(\this_ppu.M_state_q_RNISP3R6_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_4_10_LC_13_20_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_4_10_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_4_10_LC_13_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_4_10_LC_13_20_3  (
            .in0(N__21944),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21979),
            .lcout(\this_ppu.M_state_q_RNISP3R6_4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_0_10_LC_13_20_4 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_0_10_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_0_10_LC_13_20_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_0_10_LC_13_20_4  (
            .in0(N__21977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21942),
            .lcout(\this_ppu.M_state_q_RNISP3R6_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_13_20_5 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_13_20_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_13_20_5  (
            .in0(N__29809),
            .in1(N__29848),
            .in2(_gnd_net_),
            .in3(N__29821),
            .lcout(\this_ppu.N_835_0 ),
            .ltout(\this_ppu.N_835_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNINHM65_10_LC_13_20_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNINHM65_10_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNINHM65_10_LC_13_20_6 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \this_ppu.M_state_q_RNINHM65_10_LC_13_20_6  (
            .in0(N__21776),
            .in1(N__21709),
            .in2(N__21674),
            .in3(N__21608),
            .lcout(\this_ppu.N_783 ),
            .ltout(\this_ppu.N_783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNO_LC_13_20_7 .C_ON=1'b0;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNO_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNO_LC_13_20_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNO_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21671),
            .in3(N__21976),
            .lcout(\this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_13_21_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIDQQ11_LC_13_21_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIDQQ11_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(N__36546),
            .in2(_gnd_net_),
            .in3(N__36170),
            .lcout(N_92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_2_LC_13_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_2_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21662),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39360),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_0_LC_13_21_5 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_0_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_0_LC_13_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_0_LC_13_21_5  (
            .in0(N__21993),
            .in1(N__21639),
            .in2(N__21621),
            .in3(N__21476),
            .lcout(\this_ppu.N_807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_RNISP3R6_3_10_LC_13_21_6 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_RNISP3R6_3_10_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_RNISP3R6_3_10_LC_13_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_state_q_RNISP3R6_3_10_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(N__21992),
            .in2(_gnd_net_),
            .in3(N__21946),
            .lcout(\this_ppu.M_state_q_RNISP3R6_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIR9R11_LC_13_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIR9R11_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIR9R11_LC_13_22_2 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIR9R11_LC_13_22_2  (
            .in0(N__25943),
            .in1(N__25253),
            .in2(N__25304),
            .in3(N__34931),
            .lcout(N_222_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNIMU531_1_LC_13_24_4.C_ON=1'b0;
    defparam M_this_oam_address_q_RNIMU531_1_LC_13_24_4.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNIMU531_1_LC_13_24_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 M_this_oam_address_q_RNIMU531_1_LC_13_24_4 (
            .in0(N__23693),
            .in1(N__36545),
            .in2(N__23765),
            .in3(N__34926),
            .lcout(un1_M_this_oam_address_q_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_1_LC_13_26_0.C_ON=1'b0;
    defparam M_this_oam_address_q_1_LC_13_26_0.SEQ_MODE=4'b1000;
    defparam M_this_oam_address_q_1_LC_13_26_0.LUT_INIT=16'b0000011000001100;
    LogicCell40 M_this_oam_address_q_1_LC_13_26_0 (
            .in0(N__23667),
            .in1(N__23759),
            .in2(N__25216),
            .in3(N__23723),
            .lcout(M_this_oam_address_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39396),
            .ce(),
            .sr(N__38951));
    defparam M_this_data_tmp_q_esr_18_LC_13_27_3.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_18_LC_13_27_3.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_18_LC_13_27_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_18_LC_13_27_3 (
            .in0(N__37633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39402),
            .ce(N__21825),
            .sr(N__36834));
    defparam M_this_data_tmp_q_esr_1_LC_13_29_5.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_1_LC_13_29_5.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_1_LC_13_29_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_data_tmp_q_esr_1_LC_13_29_5 (
            .in0(N__37694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_data_tmp_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39409),
            .ce(N__23606),
            .sr(N__36836));
    defparam M_this_data_tmp_q_esr_19_LC_13_31_2.C_ON=1'b0;
    defparam M_this_data_tmp_q_esr_19_LC_13_31_2.SEQ_MODE=4'b1000;
    defparam M_this_data_tmp_q_esr_19_LC_13_31_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_tmp_q_esr_19_LC_13_31_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37852),
            .lcout(M_this_data_tmp_qZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39417),
            .ce(N__21849),
            .sr(N__36840));
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_14_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_3_LC_14_14_1 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_3_LC_14_14_1  (
            .in0(N__23094),
            .in1(N__22097),
            .in2(N__22134),
            .in3(N__23178),
            .lcout(this_ppu_M_screen_y_q_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39302),
            .ce(N__23059),
            .sr(N__36823));
    defparam \this_ppu.M_screen_y_q_esr_6_LC_14_14_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_6_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_6_LC_14_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_ppu.M_screen_y_q_esr_6_LC_14_14_5  (
            .in0(N__22355),
            .in1(N__22162),
            .in2(_gnd_net_),
            .in3(N__23180),
            .lcout(this_ppu_M_screen_y_q_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39302),
            .ce(N__23059),
            .sr(N__36823));
    defparam \this_ppu.M_screen_y_q_esr_7_LC_14_14_6 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_7_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_7_LC_14_14_6 .LUT_INIT=16'b0010100010100000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_7_LC_14_14_6  (
            .in0(N__23181),
            .in1(N__22356),
            .in2(N__23320),
            .in3(N__22163),
            .lcout(\this_ppu.M_screen_y_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39302),
            .ce(N__23059),
            .sr(N__36823));
    defparam \this_ppu.M_screen_y_q_esr_5_LC_14_14_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_5_LC_14_14_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_5_LC_14_14_7 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_5_LC_14_14_7  (
            .in0(N__22077),
            .in1(N__22150),
            .in2(N__22396),
            .in3(N__23179),
            .lcout(this_ppu_M_screen_y_q_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39302),
            .ce(N__23059),
            .sr(N__36823));
    defparam \this_ppu.M_screen_y_q_esr_RNIO9AV8_3_LC_14_15_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIO9AV8_3_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIO9AV8_3_LC_14_15_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIO9AV8_3_LC_14_15_2  (
            .in0(N__23140),
            .in1(N__22118),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_RNICCMV8_0_LC_14_15_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_RNICCMV8_0_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_RNICCMV8_0_LC_14_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_screen_y_q_RNICCMV8_0_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__23254),
            .in2(_gnd_net_),
            .in3(N__23139),
            .lcout(\this_ppu.M_screen_y_q_RNICCMV8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNICBI29_1_LC_14_15_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNICBI29_1_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNICBI29_1_LC_14_15_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNICBI29_1_LC_14_15_7  (
            .in0(N__23209),
            .in1(N__23253),
            .in2(_gnd_net_),
            .in3(N__23138),
            .lcout(\this_ppu.un3_M_screen_y_d_0_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIN8AV8_2_LC_14_16_0 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIN8AV8_2_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIN8AV8_2_LC_14_16_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIN8AV8_2_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__23090),
            .in2(_gnd_net_),
            .in3(N__23141),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIPAAV8_4_LC_14_16_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIPAAV8_4_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIPAAV8_4_LC_14_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIPAAV8_4_LC_14_16_1  (
            .in0(N__23142),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22084),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_2_LC_14_16_2 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_2_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_2_LC_14_16_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m68_0_a2_2_LC_14_16_2  (
            .in0(N__22043),
            .in1(N__24275),
            .in2(_gnd_net_),
            .in3(N__24059),
            .lcout(),
            .ltout(\this_ppu.m68_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_LC_14_16_3 .C_ON=1'b0;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_state_q_ns_11_0__m68_0_a2_LC_14_16_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_ppu.M_state_q_ns_11_0__m68_0_a2_LC_14_16_3  (
            .in0(N__24209),
            .in1(N__24131),
            .in2(N__22022),
            .in3(N__25010),
            .lcout(\this_ppu.M_state_q_ns_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8ES8_9_LC_14_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8ES8_9_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIM8ES8_9_LC_14_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIM8ES8_9_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__34153),
            .in2(_gnd_net_),
            .in3(N__29607),
            .lcout(M_this_ppu_vga_is_drawing),
            .ltout(M_this_ppu_vga_is_drawing_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIM7AV8_1_LC_14_16_5 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIM7AV8_1_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIM7AV8_1_LC_14_16_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIM7AV8_1_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22400),
            .in3(N__23210),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIQBAV8_5_LC_14_16_6 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIQBAV8_5_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIQBAV8_5_LC_14_16_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIQBAV8_5_LC_14_16_6  (
            .in0(N__22392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23143),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_esr_RNIRCAV8_6_LC_14_16_7 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_RNIRCAV8_6_LC_14_16_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.M_screen_y_q_esr_RNIRCAV8_6_LC_14_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_RNIRCAV8_6_LC_14_16_7  (
            .in0(N__23144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22357),
            .lcout(\this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_x_q_1_LC_14_17_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_1_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_1_LC_14_17_0 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \this_ppu.M_surface_x_q_1_LC_14_17_0  (
            .in0(N__22334),
            .in1(N__22255),
            .in2(N__22328),
            .in3(N__24865),
            .lcout(\this_ppu.M_surface_x_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39319),
            .ce(),
            .sr(N__36813));
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_14_17_1 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_14_17_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_14_17_1  (
            .in0(N__22253),
            .in1(_gnd_net_),
            .in2(N__36964),
            .in3(_gnd_net_),
            .lcout(\this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_screen_y_q_0_LC_14_17_2 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_0_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_0_LC_14_17_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \this_ppu.M_screen_y_q_0_LC_14_17_2  (
            .in0(N__23158),
            .in1(N__23241),
            .in2(N__23257),
            .in3(N__22257),
            .lcout(M_this_ppu_vram_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39319),
            .ce(),
            .sr(N__36813));
    defparam \this_ppu.M_surface_x_q_7_LC_14_17_3 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_7_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_7_LC_14_17_3 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \this_ppu.M_surface_x_q_7_LC_14_17_3  (
            .in0(N__22254),
            .in1(N__25045),
            .in2(N__22313),
            .in3(N__22304),
            .lcout(M_this_ppu_map_addr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39319),
            .ce(),
            .sr(N__36813));
    defparam \this_ppu.M_surface_x_q_4_LC_14_17_4 .C_ON=1'b0;
    defparam \this_ppu.M_surface_x_q_4_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_x_q_4_LC_14_17_4 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \this_ppu.M_surface_x_q_4_LC_14_17_4  (
            .in0(N__22295),
            .in1(N__22286),
            .in2(N__24253),
            .in3(N__22256),
            .lcout(M_this_ppu_map_addr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39319),
            .ce(),
            .sr(N__36813));
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_14_17_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_14_17_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_14_17_7  (
            .in0(N__22190),
            .in1(N__22178),
            .in2(_gnd_net_),
            .in3(N__32687),
            .lcout(M_this_ppu_spr_addr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_18_0 .C_ON=1'b1;
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__23171),
            .in2(N__23183),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_18_1 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_0_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__22751),
            .in2(N__25004),
            .in3(N__22706),
            .lcout(\this_ppu.offset_y ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_0 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_18_2 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_1_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_1_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__22703),
            .in2(N__24995),
            .in3(N__22667),
            .lcout(\this_ppu.M_surface_y_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_0 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_1 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_18_3 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_2_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_2_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__22664),
            .in2(N__24986),
            .in3(N__22625),
            .lcout(\this_ppu.M_surface_y_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_1 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_2 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_18_4 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_3_LC_14_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_3_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__22622),
            .in2(N__24977),
            .in3(N__22568),
            .lcout(M_this_ppu_map_addr_5),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_2 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_3 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_18_5 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_4_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_4_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__22565),
            .in2(N__24965),
            .in3(N__22517),
            .lcout(M_this_ppu_map_addr_6),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_3 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_4 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_18_6 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_5_LC_14_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_5_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__22514),
            .in2(N__24956),
            .in3(N__22457),
            .lcout(M_this_ppu_map_addr_7),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_4 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_5 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_18_7 .C_ON=1'b1;
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_6_LC_14_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_6_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__22454),
            .in2(N__24947),
            .in3(N__23327),
            .lcout(M_this_ppu_map_addr_8),
            .ltout(),
            .carryin(\this_ppu.un1_M_surface_y_d_cry_5 ),
            .carryout(\this_ppu.un1_M_surface_y_d_cry_6 ),
            .clk(N__39327),
            .ce(N__23058),
            .sr(N__36817));
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_19_0 .C_ON=1'b0;
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_surface_y_q_esr_7_LC_14_19_0 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \this_ppu.M_surface_y_q_esr_7_LC_14_19_0  (
            .in0(N__23177),
            .in1(N__24938),
            .in2(N__23324),
            .in3(N__23303),
            .lcout(M_this_ppu_map_addr_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39335),
            .ce(N__23051),
            .sr(N__36821));
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_19_1 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_1_LC_14_19_1 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_1_LC_14_19_1  (
            .in0(N__23255),
            .in1(N__23207),
            .in2(_gnd_net_),
            .in3(N__23175),
            .lcout(\this_ppu.M_screen_y_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39335),
            .ce(N__23051),
            .sr(N__36821));
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_19_3 .C_ON=1'b0;
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_19_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.M_screen_y_q_esr_2_LC_14_19_3 .LUT_INIT=16'b0111100000000000;
    LogicCell40 \this_ppu.M_screen_y_q_esr_2_LC_14_19_3  (
            .in0(N__23256),
            .in1(N__23208),
            .in2(N__23095),
            .in3(N__23176),
            .lcout(\this_ppu.M_screen_y_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39335),
            .ce(N__23051),
            .sr(N__36821));
    defparam CONSTANT_ONE_LUT4_LC_14_20_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_20_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_14_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIP7R11_LC_14_20_1 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIP7R11_LC_14_20_1  (
            .in0(N__25941),
            .in1(N__25248),
            .in2(N__25300),
            .in3(N__34994),
            .lcout(M_this_state_d_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_LC_14_20_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \this_start_data_delay.M_last_q_LC_14_20_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \this_start_data_delay.M_last_q_LC_14_20_2  (
            .in0(N__25249),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25291),
            .lcout(\this_start_data_delay.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39343),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_14_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_LC_14_20_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_LC_14_20_3  (
            .in0(N__25292),
            .in1(N__25937),
            .in2(_gnd_net_),
            .in3(N__25247),
            .lcout(\this_start_data_delay.N_227_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_14_20_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_14_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__23021),
            .in2(_gnd_net_),
            .in3(N__24001),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_delay_clk.M_pipe_q_4_LC_14_20_5 .C_ON=1'b0;
    defparam \this_delay_clk.M_pipe_q_4_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \this_delay_clk.M_pipe_q_4_LC_14_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_delay_clk.M_pipe_q_4_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23519),
            .lcout(M_this_delay_clk_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39343),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNILR691_2_LC_14_20_7.C_ON=1'b0;
    defparam M_this_state_q_RNILR691_2_LC_14_20_7.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNILR691_2_LC_14_20_7.LUT_INIT=16'b1110111011001100;
    LogicCell40 M_this_state_q_RNILR691_2_LC_14_20_7 (
            .in0(N__36498),
            .in1(N__36943),
            .in2(_gnd_net_),
            .in3(N__36065),
            .lcout(N_1256_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_1_LC_14_21_0.C_ON=1'b0;
    defparam M_this_data_count_q_1_LC_14_21_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_1_LC_14_21_0.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_1_LC_14_21_0 (
            .in0(N__25130),
            .in1(N__26759),
            .in2(_gnd_net_),
            .in3(N__25882),
            .lcout(M_this_data_count_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39353),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_2_LC_14_21_1.C_ON=1'b0;
    defparam M_this_data_count_q_2_LC_14_21_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_2_LC_14_21_1.LUT_INIT=16'b0100010000010001;
    LogicCell40 M_this_data_count_q_2_LC_14_21_1 (
            .in0(N__26760),
            .in1(N__25115),
            .in2(_gnd_net_),
            .in3(N__25903),
            .lcout(M_this_data_count_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39353),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_3_LC_14_21_2.C_ON=1'b0;
    defparam M_this_data_count_q_3_LC_14_21_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_3_LC_14_21_2.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_3_LC_14_21_2 (
            .in0(N__25103),
            .in1(N__26761),
            .in2(_gnd_net_),
            .in3(N__25860),
            .lcout(M_this_data_count_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39353),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_7_LC_14_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_7_LC_14_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_7_LC_14_21_3.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_7_LC_14_21_3 (
            .in0(N__26762),
            .in1(_gnd_net_),
            .in2(N__25082),
            .in3(N__26880),
            .lcout(M_this_data_count_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39353),
            .ce(N__32290),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_14_21_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_14_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__23997),
            .in2(_gnd_net_),
            .in3(N__23489),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_14_21_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_14_21_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_14_21_5  (
            .in0(N__23998),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23444),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_14_21_6 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_14_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__23999),
            .in2(_gnd_net_),
            .in3(N__23402),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_14_21_7 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_14_21_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_14_21_7  (
            .in0(N__24000),
            .in1(N__23354),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ctrl_flags_q_6_LC_14_22_0.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_6_LC_14_22_0.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_6_LC_14_22_0.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_this_ctrl_flags_q_6_LC_14_22_0 (
            .in0(N__24036),
            .in1(N__36544),
            .in2(N__37375),
            .in3(N__36032),
            .lcout(M_this_ctrl_flags_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39361),
            .ce(),
            .sr(N__36827));
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_14_25_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_14_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_14_25_2  (
            .in0(_gnd_net_),
            .in1(N__24017),
            .in2(_gnd_net_),
            .in3(N__23996),
            .lcout(\this_ppu.oam_cache.M_oam_cache_write_data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_14_26_0.C_ON=1'b0;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_14_26_0.SEQ_MODE=4'b0000;
    defparam M_this_oam_address_q_RNI24IA1_1_1_LC_14_26_0.LUT_INIT=16'b1111111100010000;
    LogicCell40 M_this_oam_address_q_RNI24IA1_1_1_LC_14_26_0 (
            .in0(N__23757),
            .in1(N__23722),
            .in2(N__23672),
            .in3(N__36934),
            .lcout(N_1248_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_2_LC_14_26_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_2_LC_14_26_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_2_LC_14_26_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_2_LC_14_26_2  (
            .in0(N__30817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25820),
            .lcout(\this_reset_cond.M_stage_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39392),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_3_LC_14_26_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_3_LC_14_26_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_3_LC_14_26_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_3_LC_14_26_4  (
            .in0(N__30818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23573),
            .lcout(\this_reset_cond.M_stage_qZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39392),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK6R81_1_LC_15_15_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_1_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_1_LC_15_15_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK6R81_1_LC_15_15_4  (
            .in0(N__36539),
            .in1(N__35633),
            .in2(_gnd_net_),
            .in3(N__38277),
            .lcout(M_this_spr_ram_write_en_0_i_1_0),
            .ltout(M_this_spr_ram_write_en_0_i_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_15_15_5 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_6_0_wclke_3_LC_15_15_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_spr_ram.mem_mem_6_0_wclke_3_LC_15_15_5  (
            .in0(N__32000),
            .in1(N__32204),
            .in2(N__23567),
            .in3(N__32102),
            .lcout(\this_spr_ram.mem_WE_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_15_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_15_16_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_15_16_1  (
            .in0(N__31226),
            .in1(N__26535),
            .in2(N__31354),
            .in3(N__26659),
            .lcout(\this_vga_signals.M_vcounter_d7lt8_0 ),
            .ltout(\this_vga_signals.M_vcounter_d7lt8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_16_2 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_16_2  (
            .in0(N__26393),
            .in1(N__33940),
            .in2(N__24932),
            .in3(N__35271),
            .lcout(\this_vga_signals.M_vcounter_d8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_15_17_0 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_0_c_inv_LC_15_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.offset_x_cry_0_c_inv_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__24884),
            .in2(N__24929),
            .in3(N__26554),
            .lcout(\this_ppu.M_oam_cache_read_data_i_8 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\this_ppu.offset_x_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_15_17_1 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_15_17_1 .LUT_INIT=16'b1110000110110100;
    LogicCell40 \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_15_17_1  (
            .in0(N__32680),
            .in1(N__24878),
            .in2(N__24866),
            .in3(N__24590),
            .lcout(M_this_ppu_spr_addr_1),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_0 ),
            .carryout(\this_ppu.offset_x_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_15_17_2 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_15_17_2 .LUT_INIT=16'b1110000110110100;
    LogicCell40 \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_15_17_2  (
            .in0(N__32694),
            .in1(N__24587),
            .in2(N__24578),
            .in3(N__24332),
            .lcout(M_this_ppu_spr_addr_2),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_1 ),
            .carryout(\this_ppu.offset_x_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_2_c_RNI0QAP_LC_15_17_3 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_2_c_RNI0QAP_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_2_c_RNI0QAP_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_2_c_RNI0QAP_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__26363),
            .in2(N__24328),
            .in3(N__24269),
            .lcout(\this_ppu.offset_x_3 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_2 ),
            .carryout(\this_ppu.offset_x_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_15_17_4 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__26591),
            .in2(N__24252),
            .in3(N__24203),
            .lcout(\this_ppu.offset_x_4 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_3 ),
            .carryout(\this_ppu.offset_x_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_15_17_5 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_4_c_RNI62DP_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_4_c_RNI62DP_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__24200),
            .in2(N__24181),
            .in3(N__24125),
            .lcout(\this_ppu.offset_x_5 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_4 ),
            .carryout(\this_ppu.offset_x_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_15_17_6 .C_ON=1'b1;
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_5_c_RNI96EP_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \this_ppu.offset_x_cry_5_c_RNI96EP_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__24122),
            .in2(N__24103),
            .in3(N__24053),
            .lcout(\this_ppu.offset_x_6 ),
            .ltout(),
            .carryin(\this_ppu.offset_x_cry_5 ),
            .carryout(\this_ppu.offset_x_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_15_17_7 .C_ON=1'b0;
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \this_ppu.offset_x_cry_6_c_RNICAFP_LC_15_17_7 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \this_ppu.offset_x_cry_6_c_RNICAFP_LC_15_17_7  (
            .in0(N__25044),
            .in1(_gnd_net_),
            .in2(N__25025),
            .in3(N__25013),
            .lcout(\this_ppu.offset_x_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_scroll_q_esr_0_LC_15_18_0.C_ON=1'b0;
    defparam M_this_scroll_q_esr_0_LC_15_18_0.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_0_LC_15_18_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_0_LC_15_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38128),
            .lcout(M_this_scroll_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_1_LC_15_18_1.C_ON=1'b0;
    defparam M_this_scroll_q_esr_1_LC_15_18_1.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_1_LC_15_18_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_1_LC_15_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37759),
            .lcout(M_this_scroll_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_2_LC_15_18_2.C_ON=1'b0;
    defparam M_this_scroll_q_esr_2_LC_15_18_2.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_2_LC_15_18_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_2_LC_15_18_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37628),
            .lcout(M_this_scroll_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_3_LC_15_18_3.C_ON=1'b0;
    defparam M_this_scroll_q_esr_3_LC_15_18_3.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_3_LC_15_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_3_LC_15_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37879),
            .lcout(M_this_scroll_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_4_LC_15_18_4.C_ON=1'b0;
    defparam M_this_scroll_q_esr_4_LC_15_18_4.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_4_LC_15_18_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_4_LC_15_18_4 (
            .in0(N__37520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_5_LC_15_18_5.C_ON=1'b0;
    defparam M_this_scroll_q_esr_5_LC_15_18_5.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_5_LC_15_18_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_5_LC_15_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38890),
            .lcout(M_this_scroll_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_6_LC_15_18_6.C_ON=1'b0;
    defparam M_this_scroll_q_esr_6_LC_15_18_6.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_6_LC_15_18_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_scroll_q_esr_6_LC_15_18_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37351),
            .lcout(M_this_scroll_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_scroll_q_esr_7_LC_15_18_7.C_ON=1'b0;
    defparam M_this_scroll_q_esr_7_LC_15_18_7.SEQ_MODE=4'b1000;
    defparam M_this_scroll_q_esr_7_LC_15_18_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 M_this_scroll_q_esr_7_LC_15_18_7 (
            .in0(N__38759),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(M_this_scroll_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39320),
            .ce(N__35522),
            .sr(N__36814));
    defparam M_this_data_count_q_cry_c_0_LC_15_19_0.C_ON=1'b1;
    defparam M_this_data_count_q_cry_c_0_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_c_0_LC_15_19_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 M_this_data_count_q_cry_c_0_LC_15_19_0 (
            .in0(_gnd_net_),
            .in1(N__25838),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(M_this_data_count_q_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_15_19_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_0_THRU_LUT4_0_LC_15_19_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_0_THRU_LUT4_0_LC_15_19_1 (
            .in0(_gnd_net_),
            .in1(N__25883),
            .in2(N__25402),
            .in3(N__25118),
            .lcout(M_this_data_count_q_cry_0_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_0),
            .carryout(M_this_data_count_q_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_15_19_2.C_ON=1'b1;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_1_THRU_LUT4_0_LC_15_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_1_THRU_LUT4_0_LC_15_19_2 (
            .in0(_gnd_net_),
            .in1(N__25370),
            .in2(N__25907),
            .in3(N__25106),
            .lcout(M_this_data_count_q_cry_1_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_1),
            .carryout(M_this_data_count_q_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_15_19_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_2_THRU_LUT4_0_LC_15_19_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_2_THRU_LUT4_0_LC_15_19_3 (
            .in0(_gnd_net_),
            .in1(N__25862),
            .in2(N__25403),
            .in3(N__25094),
            .lcout(M_this_data_count_q_cry_2_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_2),
            .carryout(M_this_data_count_q_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_15_19_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_3_THRU_LUT4_0_LC_15_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_3_THRU_LUT4_0_LC_15_19_4 (
            .in0(_gnd_net_),
            .in1(N__25374),
            .in2(N__26021),
            .in3(N__25091),
            .lcout(M_this_data_count_q_cry_3_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_3),
            .carryout(M_this_data_count_q_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_15_19_5.C_ON=1'b1;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_4_THRU_LUT4_0_LC_15_19_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_4_THRU_LUT4_0_LC_15_19_5 (
            .in0(_gnd_net_),
            .in1(N__25988),
            .in2(N__25404),
            .in3(N__25088),
            .lcout(M_this_data_count_q_cry_4_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_4),
            .carryout(M_this_data_count_q_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_15_19_6.C_ON=1'b1;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_15_19_6.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_5_THRU_LUT4_0_LC_15_19_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_5_THRU_LUT4_0_LC_15_19_6 (
            .in0(_gnd_net_),
            .in1(N__25378),
            .in2(N__26714),
            .in3(N__25085),
            .lcout(M_this_data_count_q_cry_5_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_5),
            .carryout(M_this_data_count_q_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_15_19_7.C_ON=1'b1;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_6_THRU_LUT4_0_LC_15_19_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_6_THRU_LUT4_0_LC_15_19_7 (
            .in0(_gnd_net_),
            .in1(N__26882),
            .in2(N__25405),
            .in3(N__25070),
            .lcout(M_this_data_count_q_cry_6_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_6),
            .carryout(M_this_data_count_q_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_8_LC_15_20_0.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_8_LC_15_20_0.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_8_LC_15_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_8_LC_15_20_0 (
            .in0(_gnd_net_),
            .in1(N__25142),
            .in2(N__25400),
            .in3(N__25067),
            .lcout(M_this_data_count_q_s_8),
            .ltout(),
            .carryin(bfn_15_20_0_),
            .carryout(M_this_data_count_q_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_15_20_1.C_ON=1'b1;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_8_THRU_LUT4_0_LC_15_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_8_THRU_LUT4_0_LC_15_20_1 (
            .in0(_gnd_net_),
            .in1(N__25366),
            .in2(N__25964),
            .in3(N__25814),
            .lcout(M_this_data_count_q_cry_8_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_8),
            .carryout(M_this_data_count_q_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_10_LC_15_20_2.C_ON=1'b1;
    defparam M_this_data_count_q_RNO_0_10_LC_15_20_2.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_10_LC_15_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 M_this_data_count_q_RNO_0_10_LC_15_20_2 (
            .in0(_gnd_net_),
            .in1(N__26792),
            .in2(N__25399),
            .in3(N__25811),
            .lcout(M_this_data_count_q_s_10),
            .ltout(),
            .carryin(M_this_data_count_q_cry_9),
            .carryout(M_this_data_count_q_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_15_20_3.C_ON=1'b1;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_15_20_3.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_10_THRU_LUT4_0_LC_15_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_10_THRU_LUT4_0_LC_15_20_3 (
            .in0(_gnd_net_),
            .in1(N__25362),
            .in2(N__26825),
            .in3(N__25808),
            .lcout(M_this_data_count_q_cry_10_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_10),
            .carryout(M_this_data_count_q_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_15_20_4.C_ON=1'b1;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_cry_11_THRU_LUT4_0_LC_15_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 M_this_data_count_q_cry_11_THRU_LUT4_0_LC_15_20_4 (
            .in0(_gnd_net_),
            .in1(N__26840),
            .in2(N__25401),
            .in3(N__25310),
            .lcout(M_this_data_count_q_cry_11_THRU_CO),
            .ltout(),
            .carryin(M_this_data_count_q_cry_11),
            .carryout(M_this_data_count_q_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_RNO_0_13_LC_15_20_5.C_ON=1'b0;
    defparam M_this_data_count_q_RNO_0_13_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam M_this_data_count_q_RNO_0_13_LC_15_20_5.LUT_INIT=16'b1100110000110011;
    LogicCell40 M_this_data_count_q_RNO_0_13_LC_15_20_5 (
            .in0(_gnd_net_),
            .in1(N__26806),
            .in2(_gnd_net_),
            .in3(N__25307),
            .lcout(M_this_data_count_q_s_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_15_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_15_20_6 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_15_20_6  (
            .in0(N__25296),
            .in1(N__25936),
            .in2(_gnd_net_),
            .in3(N__25246),
            .lcout(N_220_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_9_LC_15_20_7.C_ON=1'b0;
    defparam M_this_state_q_9_LC_15_20_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_9_LC_15_20_7.LUT_INIT=16'b0010001000000000;
    LogicCell40 M_this_state_q_9_LC_15_20_7 (
            .in0(N__36502),
            .in1(N__36957),
            .in2(_gnd_net_),
            .in3(N__35621),
            .lcout(M_this_state_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39336),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_8_LC_15_21_0.C_ON=1'b0;
    defparam M_this_data_count_q_8_LC_15_21_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_8_LC_15_21_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 M_this_data_count_q_8_LC_15_21_0 (
            .in0(N__36949),
            .in1(N__25226),
            .in2(N__25211),
            .in3(N__26753),
            .lcout(M_this_data_count_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39344),
            .ce(N__32294),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_7_11_LC_15_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_7_11_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_7_11_LC_15_21_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_7_11_LC_15_21_1  (
            .in0(N__25141),
            .in1(N__25983),
            .in2(N__25963),
            .in3(N__26013),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_4_LC_15_21_2.C_ON=1'b0;
    defparam M_this_data_count_q_4_LC_15_21_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_4_LC_15_21_2.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_4_LC_15_21_2 (
            .in0(N__26014),
            .in1(N__26033),
            .in2(_gnd_net_),
            .in3(N__26750),
            .lcout(M_this_data_count_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39344),
            .ce(N__32294),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_5_LC_15_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_5_LC_15_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_5_LC_15_21_3.LUT_INIT=16'b0101000000000101;
    LogicCell40 M_this_data_count_q_5_LC_15_21_3 (
            .in0(N__26751),
            .in1(_gnd_net_),
            .in2(N__26000),
            .in3(N__25984),
            .lcout(M_this_data_count_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39344),
            .ce(N__32294),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_9_LC_15_21_4.C_ON=1'b0;
    defparam M_this_data_count_q_9_LC_15_21_4.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_9_LC_15_21_4.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_9_LC_15_21_4 (
            .in0(N__25970),
            .in1(N__26752),
            .in2(_gnd_net_),
            .in3(N__25959),
            .lcout(M_this_data_count_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39344),
            .ce(N__32294),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI30CP2_LC_15_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI30CP2_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI30CP2_LC_15_21_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \this_start_data_delay.M_last_q_RNI30CP2_LC_15_21_5  (
            .in0(N__38308),
            .in1(N__25942),
            .in2(_gnd_net_),
            .in3(N__36948),
            .lcout(N_685_i),
            .ltout(N_685_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_0_LC_15_21_6.C_ON=1'b0;
    defparam M_this_data_count_q_0_LC_15_21_6.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_0_LC_15_21_6.LUT_INIT=16'b0000100100001001;
    LogicCell40 M_this_data_count_q_0_LC_15_21_6 (
            .in0(N__25834),
            .in1(_gnd_net_),
            .in2(N__25910),
            .in3(_gnd_net_),
            .lcout(M_this_data_count_qZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39344),
            .ce(N__32294),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_9_11_LC_15_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_9_11_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_9_11_LC_15_21_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_9_11_LC_15_21_7  (
            .in0(N__25899),
            .in1(N__25878),
            .in2(N__25861),
            .in3(N__25833),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_5_LC_15_25_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_5_LC_15_25_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_5_LC_15_25_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \this_reset_cond.M_stage_q_5_LC_15_25_2  (
            .in0(_gnd_net_),
            .in1(N__26336),
            .in2(_gnd_net_),
            .in3(N__30801),
            .lcout(\this_reset_cond.M_stage_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39376),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_1_LC_15_26_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_1_LC_15_26_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_1_LC_15_26_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_1_LC_15_26_0  (
            .in0(N__30815),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26330),
            .lcout(\this_reset_cond.M_stage_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39384),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_4_LC_15_26_1 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_4_LC_15_26_1 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_4_LC_15_26_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_4_LC_15_26_1  (
            .in0(_gnd_net_),
            .in1(N__30816),
            .in2(_gnd_net_),
            .in3(N__26342),
            .lcout(\this_reset_cond.M_stage_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39384),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_0_LC_15_26_2 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_0_LC_15_26_2 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_0_LC_15_26_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \this_reset_cond.M_stage_q_0_LC_15_26_2  (
            .in0(N__30814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_reset_cond.M_stage_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39384),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_16_13_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_16_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_16_13_4  (
            .in0(N__26051),
            .in1(N__26324),
            .in2(_gnd_net_),
            .in3(N__32701),
            .lcout(M_this_ppu_spr_addr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_0_LC_16_13_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_0_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_0_LC_16_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_0_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26066),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39288),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_0_LC_16_15_0 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_0_LC_16_15_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_0_LC_16_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_0_LC_16_15_0  (
            .in0(N__29770),
            .in1(N__26536),
            .in2(N__28616),
            .in3(N__28611),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .clk(N__39296),
            .ce(),
            .sr(N__34426));
    defparam \this_vga_signals.M_vcounter_q_1_LC_16_15_1 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_1_LC_16_15_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_1_LC_16_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_1_LC_16_15_1  (
            .in0(N__29772),
            .in1(N__26666),
            .in2(_gnd_net_),
            .in3(N__26045),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_1 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_0 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .clk(N__39296),
            .ce(),
            .sr(N__34426));
    defparam \this_vga_signals.M_vcounter_q_2_LC_16_15_2 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_2_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_2_LC_16_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_2_LC_16_15_2  (
            .in0(N__29771),
            .in1(N__31260),
            .in2(_gnd_net_),
            .in3(N__26042),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_2 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_1 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .clk(N__39296),
            .ce(),
            .sr(N__34426));
    defparam \this_vga_signals.M_vcounter_q_3_LC_16_15_3 .C_ON=1'b1;
    defparam \this_vga_signals.M_vcounter_q_3_LC_16_15_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_3_LC_16_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_3_LC_16_15_3  (
            .in0(N__29773),
            .in1(N__31352),
            .in2(_gnd_net_),
            .in3(N__26039),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_3 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_2 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .clk(N__39296),
            .ce(),
            .sr(N__34426));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_16_15_4 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_16_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__33941),
            .in2(_gnd_net_),
            .in3(N__26036),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_3 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_16_15_5 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_16_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__33184),
            .in2(_gnd_net_),
            .in3(N__26408),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_4 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_16_15_6 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_16_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__34061),
            .in2(_gnd_net_),
            .in3(N__26405),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_5 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_16_15_7 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_16_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__34754),
            .in2(_gnd_net_),
            .in3(N__26402),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0 ),
            .ltout(),
            .carryin(\this_vga_signals.un1_M_vcounter_q_cry_6 ),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_16_16_0 .C_ON=1'b1;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_16_16_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34655),
            .in3(N__26399),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\this_vga_signals.un1_M_vcounter_q_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_16_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_16_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__35272),
            .in2(_gnd_net_),
            .in3(N__26396),
            .lcout(\this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNILL3J1_1_LC_16_16_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNILL3J1_1_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNILL3J1_1_LC_16_16_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNILL3J1_1_LC_16_16_4  (
            .in0(N__31353),
            .in1(N__26667),
            .in2(N__34753),
            .in3(N__33925),
            .lcout(\this_vga_signals.m43_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_16_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_16_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_16_16_5  (
            .in0(N__34060),
            .in1(N__34651),
            .in2(N__33183),
            .in3(N__34745),
            .lcout(\this_vga_signals.M_vcounter_d7lto9_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPIAB9_9_LC_16_16_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPIAB9_9_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIPIAB9_9_LC_16_16_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIPIAB9_9_LC_16_16_6  (
            .in0(N__28538),
            .in1(N__34154),
            .in2(_gnd_net_),
            .in3(N__29598),
            .lcout(port_nmib_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_16_17_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI72M7_11_LC_16_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI72M7_11_LC_16_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26609),
            .lcout(\this_ppu.M_oam_cache_read_data_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_11_LC_16_17_2 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_11_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_11_LC_16_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_11_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26357),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39305),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_16_17_5 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI83M7_12_LC_16_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI83M7_12_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26603),
            .lcout(\this_ppu.M_oam_cache_read_data_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_8_LC_16_18_4 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_8_LC_16_18_4 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_8_LC_16_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_ppu.oam_cache.read_data_8_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26585),
            .lcout(\this_ppu.M_oam_cache_read_data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39308),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_N_2L1_LC_16_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_2L1_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_2L1_LC_16_18_6 .LUT_INIT=16'b0010001001000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_N_2L1_LC_16_18_6  (
            .in0(N__30488),
            .in1(N__31523),
            .in2(_gnd_net_),
            .in3(N__30581),
            .lcout(\this_vga_signals.g0_41_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_LC_16_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_LC_16_19_0 .LUT_INIT=16'b1011100001000111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_LC_16_19_0  (
            .in0(N__30417),
            .in1(N__29966),
            .in2(N__30287),
            .in3(N__26504),
            .lcout(),
            .ltout(\this_vga_signals.N_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_16_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_15_LC_16_19_1 .LUT_INIT=16'b1110010110000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_15_LC_16_19_1  (
            .in0(N__26669),
            .in1(N__26543),
            .in2(N__26519),
            .in3(N__31187),
            .lcout(\this_vga_signals.mult1_un82_sum_c3_0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_LC_16_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_LC_16_19_2 .LUT_INIT=16'b0101000010101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_N_4L5_LC_16_19_2  (
            .in0(N__31405),
            .in1(_gnd_net_),
            .in2(N__30419),
            .in3(N__30002),
            .lcout(),
            .ltout(\this_vga_signals.g0_41_N_4L5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_1_LC_16_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_1_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_1_LC_16_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_1_LC_16_19_3  (
            .in0(N__31286),
            .in1(N__26516),
            .in2(N__26507),
            .in3(N__29891),
            .lcout(\this_vga_signals.g0_41_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNI8D7RUG1_2_LC_16_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNI8D7RUG1_2_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNI8D7RUG1_2_LC_16_19_4 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNI8D7RUG1_2_LC_16_19_4  (
            .in0(N__30047),
            .in1(N__29912),
            .in2(N__26498),
            .in3(N__26432),
            .lcout(M_this_vga_signals_address_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIVIOMG4_2_LC_16_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIVIOMG4_2_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIVIOMG4_2_LC_16_19_5 .LUT_INIT=16'b1000110000111011;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIVIOMG4_2_LC_16_19_5  (
            .in0(N__31287),
            .in1(N__29996),
            .in2(N__26624),
            .in3(N__31406),
            .lcout(\this_vga_signals.mult1_un68_sum_c3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_4_LC_16_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_4_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_4_LC_16_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x2_4_LC_16_20_0  (
            .in0(N__30501),
            .in1(N__30223),
            .in2(N__30017),
            .in3(N__30590),
            .lcout(\this_vga_signals.g0_i_x2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_16_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_LC_16_20_1 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_LC_16_20_1  (
            .in0(N__31739),
            .in1(N__31094),
            .in2(N__30230),
            .in3(N__29960),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_16_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_LC_16_20_2 .LUT_INIT=16'b1101101110111101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_LC_16_20_2  (
            .in0(N__26668),
            .in1(N__31288),
            .in2(N__26636),
            .in3(N__26633),
            .lcout(\this_vga_signals.if_m5_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_16_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBOQ11_LC_16_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBOQ11_LC_16_20_3  (
            .in0(N__36494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38171),
            .lcout(N_241_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_16_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_18_LC_16_20_4 .LUT_INIT=16'b0000010101000010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_18_LC_16_20_4  (
            .in0(N__33608),
            .in1(N__33410),
            .in2(N__33185),
            .in3(N__30623),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_16_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_3_LC_16_20_5 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_3_LC_16_20_5  (
            .in0(N__33938),
            .in1(_gnd_net_),
            .in2(N__26627),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2UNG73_4_LC_16_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2UNG73_4_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI2UNG73_4_LC_16_20_6 .LUT_INIT=16'b1010010101100101;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI2UNG73_4_LC_16_20_6  (
            .in0(N__29906),
            .in1(N__31738),
            .in2(N__33209),
            .in3(N__30222),
            .lcout(\this_vga_signals.N_17_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g2_1_2_LC_16_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g2_1_2_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g2_1_2_LC_16_20_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g2_1_2_LC_16_20_7  (
            .in0(N__33409),
            .in1(N__34045),
            .in2(N__33944),
            .in3(N__33607),
            .lcout(\this_vga_signals.g2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_10_LC_16_21_0.C_ON=1'b0;
    defparam M_this_data_count_q_10_LC_16_21_0.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_10_LC_16_21_0.LUT_INIT=16'b0100010011100100;
    LogicCell40 M_this_data_count_q_10_LC_16_21_0 (
            .in0(N__26757),
            .in1(N__26615),
            .in2(N__39530),
            .in3(N__36961),
            .lcout(M_this_data_count_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39330),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_12_LC_16_21_1.C_ON=1'b0;
    defparam M_this_data_count_q_12_LC_16_21_1.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_12_LC_16_21_1.LUT_INIT=16'b0010001000010001;
    LogicCell40 M_this_data_count_q_12_LC_16_21_1 (
            .in0(N__26900),
            .in1(N__26755),
            .in2(_gnd_net_),
            .in3(N__26839),
            .lcout(M_this_data_count_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39330),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_13_LC_16_21_2.C_ON=1'b0;
    defparam M_this_data_count_q_13_LC_16_21_2.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_13_LC_16_21_2.LUT_INIT=16'b0100010011100100;
    LogicCell40 M_this_data_count_q_13_LC_16_21_2 (
            .in0(N__26758),
            .in1(N__26894),
            .in2(N__35777),
            .in3(N__36962),
            .lcout(M_this_data_count_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39330),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_11_LC_16_21_3.C_ON=1'b0;
    defparam M_this_data_count_q_11_LC_16_21_3.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_11_LC_16_21_3.LUT_INIT=16'b0000000010011001;
    LogicCell40 M_this_data_count_q_11_LC_16_21_3 (
            .in0(N__26821),
            .in1(N__26888),
            .in2(_gnd_net_),
            .in3(N__26754),
            .lcout(M_this_data_count_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39330),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_6_11_LC_16_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_6_11_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_6_11_LC_16_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_6_11_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__26881),
            .in2(_gnd_net_),
            .in3(N__26703),
            .lcout(),
            .ltout(\this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_11_LC_16_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_11_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_11_LC_16_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_11_LC_16_21_5  (
            .in0(N__26858),
            .in1(N__26780),
            .in2(N__26849),
            .in3(N__26846),
            .lcout(N_930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_8_11_LC_16_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_8_11_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_q_srsts_i_a2_0_8_11_LC_16_21_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_this_state_q_srsts_i_a2_0_8_11_LC_16_21_6  (
            .in0(N__26838),
            .in1(N__26820),
            .in2(N__26807),
            .in3(N__26791),
            .lcout(\this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_data_count_q_6_LC_16_21_7.C_ON=1'b0;
    defparam M_this_data_count_q_6_LC_16_21_7.SEQ_MODE=4'b1000;
    defparam M_this_data_count_q_6_LC_16_21_7.LUT_INIT=16'b0000000010100101;
    LogicCell40 M_this_data_count_q_6_LC_16_21_7 (
            .in0(N__26704),
            .in1(_gnd_net_),
            .in2(N__26774),
            .in3(N__26756),
            .lcout(M_this_data_count_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39330),
            .ce(N__32286),
            .sr(_gnd_net_));
    defparam M_this_ctrl_flags_q_5_LC_16_22_5.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_5_LC_16_22_5.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_5_LC_16_22_5.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_this_ctrl_flags_q_5_LC_16_22_5 (
            .in0(N__26683),
            .in1(N__36551),
            .in2(N__38909),
            .in3(N__36034),
            .lcout(M_this_ctrl_flags_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39338),
            .ce(),
            .sr(N__36824));
    defparam M_this_ctrl_flags_q_7_LC_16_22_6.C_ON=1'b0;
    defparam M_this_ctrl_flags_q_7_LC_16_22_6.SEQ_MODE=4'b1000;
    defparam M_this_ctrl_flags_q_7_LC_16_22_6.LUT_INIT=16'b1101100011110000;
    LogicCell40 M_this_ctrl_flags_q_7_LC_16_22_6 (
            .in0(N__36033),
            .in1(N__38761),
            .in2(N__28534),
            .in3(N__36552),
            .lcout(M_this_ctrl_flags_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39338),
            .ce(),
            .sr(N__36824));
    defparam \this_reset_cond.M_stage_q_6_LC_16_23_5 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_6_LC_16_23_5 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_6_LC_16_23_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_6_LC_16_23_5  (
            .in0(N__30781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28517),
            .lcout(\this_reset_cond.M_stage_qZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39349),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_spr_address_q_0_LC_17_12_0.C_ON=1'b1;
    defparam M_this_spr_address_q_0_LC_17_12_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_0_LC_17_12_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_0_LC_17_12_0 (
            .in0(N__35806),
            .in1(N__28302),
            .in2(N__28673),
            .in3(N__28672),
            .lcout(M_this_spr_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(un1_M_this_spr_address_q_cry_0),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_1_LC_17_12_1.C_ON=1'b1;
    defparam M_this_spr_address_q_1_LC_17_12_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_1_LC_17_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_1_LC_17_12_1 (
            .in0(N__35810),
            .in1(N__28073),
            .in2(_gnd_net_),
            .in3(N__28058),
            .lcout(M_this_spr_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_0),
            .carryout(un1_M_this_spr_address_q_cry_1),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_2_LC_17_12_2.C_ON=1'b1;
    defparam M_this_spr_address_q_2_LC_17_12_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_2_LC_17_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_2_LC_17_12_2 (
            .in0(N__35807),
            .in1(N__27859),
            .in2(_gnd_net_),
            .in3(N__27809),
            .lcout(M_this_spr_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_1),
            .carryout(un1_M_this_spr_address_q_cry_2),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_3_LC_17_12_3.C_ON=1'b1;
    defparam M_this_spr_address_q_3_LC_17_12_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_3_LC_17_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_3_LC_17_12_3 (
            .in0(N__35811),
            .in1(N__27600),
            .in2(_gnd_net_),
            .in3(N__27569),
            .lcout(M_this_spr_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_2),
            .carryout(un1_M_this_spr_address_q_cry_3),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_4_LC_17_12_4.C_ON=1'b1;
    defparam M_this_spr_address_q_4_LC_17_12_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_4_LC_17_12_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_4_LC_17_12_4 (
            .in0(N__35808),
            .in1(N__27371),
            .in2(_gnd_net_),
            .in3(N__27347),
            .lcout(M_this_spr_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_3),
            .carryout(un1_M_this_spr_address_q_cry_4),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_5_LC_17_12_5.C_ON=1'b1;
    defparam M_this_spr_address_q_5_LC_17_12_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_5_LC_17_12_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_5_LC_17_12_5 (
            .in0(N__35812),
            .in1(N__27182),
            .in2(_gnd_net_),
            .in3(N__27140),
            .lcout(M_this_spr_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_4),
            .carryout(un1_M_this_spr_address_q_cry_5),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_6_LC_17_12_6.C_ON=1'b1;
    defparam M_this_spr_address_q_6_LC_17_12_6.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_6_LC_17_12_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_6_LC_17_12_6 (
            .in0(N__35809),
            .in1(N__26928),
            .in2(_gnd_net_),
            .in3(N__26903),
            .lcout(M_this_spr_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_5),
            .carryout(un1_M_this_spr_address_q_cry_6),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_7_LC_17_12_7.C_ON=1'b1;
    defparam M_this_spr_address_q_7_LC_17_12_7.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_7_LC_17_12_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_7_LC_17_12_7 (
            .in0(N__35813),
            .in1(N__29401),
            .in2(_gnd_net_),
            .in3(N__29357),
            .lcout(M_this_spr_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_6),
            .carryout(un1_M_this_spr_address_q_cry_7),
            .clk(N__39290),
            .ce(),
            .sr(N__38961));
    defparam M_this_spr_address_q_8_LC_17_13_0.C_ON=1'b1;
    defparam M_this_spr_address_q_8_LC_17_13_0.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_8_LC_17_13_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_8_LC_17_13_0 (
            .in0(N__35783),
            .in1(N__29192),
            .in2(_gnd_net_),
            .in3(N__29150),
            .lcout(M_this_spr_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(un1_M_this_spr_address_q_cry_8),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam M_this_spr_address_q_9_LC_17_13_1.C_ON=1'b1;
    defparam M_this_spr_address_q_9_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_9_LC_17_13_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_9_LC_17_13_1 (
            .in0(N__35786),
            .in1(N__28959),
            .in2(_gnd_net_),
            .in3(N__28916),
            .lcout(M_this_spr_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_8),
            .carryout(un1_M_this_spr_address_q_cry_9),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam M_this_spr_address_q_10_LC_17_13_2.C_ON=1'b1;
    defparam M_this_spr_address_q_10_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_10_LC_17_13_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_10_LC_17_13_2 (
            .in0(N__35781),
            .in1(N__28722),
            .in2(_gnd_net_),
            .in3(N__28685),
            .lcout(M_this_spr_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_9),
            .carryout(un1_M_this_spr_address_q_cry_10),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam M_this_spr_address_q_11_LC_17_13_3.C_ON=1'b1;
    defparam M_this_spr_address_q_11_LC_17_13_3.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_11_LC_17_13_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_11_LC_17_13_3 (
            .in0(N__35785),
            .in1(N__32080),
            .in2(_gnd_net_),
            .in3(N__28682),
            .lcout(M_this_spr_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_10),
            .carryout(un1_M_this_spr_address_q_cry_11),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam M_this_spr_address_q_12_LC_17_13_4.C_ON=1'b1;
    defparam M_this_spr_address_q_12_LC_17_13_4.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_12_LC_17_13_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_spr_address_q_12_LC_17_13_4 (
            .in0(N__35782),
            .in1(N__32176),
            .in2(_gnd_net_),
            .in3(N__28679),
            .lcout(M_this_spr_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_spr_address_q_cry_11),
            .carryout(un1_M_this_spr_address_q_cry_12),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam M_this_spr_address_q_13_LC_17_13_5.C_ON=1'b0;
    defparam M_this_spr_address_q_13_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam M_this_spr_address_q_13_LC_17_13_5.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_spr_address_q_13_LC_17_13_5 (
            .in0(N__31972),
            .in1(N__35784),
            .in2(_gnd_net_),
            .in3(N__28676),
            .lcout(M_this_spr_address_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39293),
            .ce(),
            .sr(N__38958));
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_17_15_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_LC_17_15_1 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK6R81_LC_17_15_1  (
            .in0(N__38282),
            .in1(N__36567),
            .in2(_gnd_net_),
            .in3(N__35629),
            .lcout(M_this_spr_ram_write_en_0_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNINK957_9_LC_17_15_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINK957_9_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNINK957_9_LC_17_15_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNINK957_9_LC_17_15_6  (
            .in0(N__28647),
            .in1(N__28610),
            .in2(_gnd_net_),
            .in3(N__29766),
            .lcout(\this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_2_LC_17_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_2_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIOLTE3_2_LC_17_16_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIOLTE3_2_LC_17_16_1  (
            .in0(N__29885),
            .in1(N__30086),
            .in2(N__31272),
            .in3(N__34041),
            .lcout(this_vga_signals_vsync_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.line_clk.M_last_q_LC_17_16_3 .C_ON=1'b0;
    defparam \this_ppu.line_clk.M_last_q_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.line_clk.M_last_q_LC_17_16_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_ppu.line_clk.M_last_q_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__29855),
            .in2(_gnd_net_),
            .in3(N__29828),
            .lcout(\this_ppu.line_clk.M_last_qZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39307),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNICF6E7_9_LC_17_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICF6E7_9_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNICF6E7_9_LC_17_16_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNICF6E7_9_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__29790),
            .in2(_gnd_net_),
            .in3(N__29650),
            .lcout(\this_vga_signals.N_933_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_36_LC_17_17_2 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_36_LC_17_17_2  (
            .in0(N__33123),
            .in1(N__33000),
            .in2(_gnd_net_),
            .in3(N__32935),
            .lcout(\this_vga_signals.N_10_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_1_LC_17_17_3 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_1_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \this_ppu.oam_cache.read_data_1_LC_17_17_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_1_LC_17_17_3  (
            .in0(N__29636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_ppu.oam_cache.M_oam_cache_read_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39313),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB4G42_9_LC_17_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB4G42_9_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIB4G42_9_LC_17_17_6 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIB4G42_9_LC_17_17_6  (
            .in0(N__34633),
            .in1(N__35257),
            .in2(N__30080),
            .in3(N__34732),
            .lcout(),
            .ltout(\this_vga_signals.vvisibility_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_9_LC_17_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_9_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_9_LC_17_17_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_9_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29621),
            .in3(N__31159),
            .lcout(\this_vga_signals.vvisibility ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_17_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_4_LC_17_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_4_LC_17_18_3  (
            .in0(N__33687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39321),
            .ce(N__34484),
            .sr(N__34427));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_1_LC_17_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_1_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_1_LC_17_18_4 .LUT_INIT=16'b0000001001011111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_0_1_LC_17_18_4  (
            .in0(N__33907),
            .in1(N__33126),
            .in2(N__34065),
            .in3(N__33610),
            .lcout(\this_vga_signals.g0_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_x2_0_LC_17_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_x2_0_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_x2_0_LC_17_18_5 .LUT_INIT=16'b0101010110011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_x2_0_LC_17_18_5  (
            .in0(N__33127),
            .in1(N__33002),
            .in2(_gnd_net_),
            .in3(N__32934),
            .lcout(),
            .ltout(\this_vga_signals.N_10_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_LC_17_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_0_LC_17_18_6 .LUT_INIT=16'b1000100001000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_0_LC_17_18_6  (
            .in0(N__29954),
            .in1(N__33408),
            .in2(N__29948),
            .in3(N__33611),
            .lcout(),
            .ltout(\this_vga_signals.g0_0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_6_LC_17_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_6_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_6_LC_17_18_7 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_6_LC_17_18_7  (
            .in0(N__29945),
            .in1(N__29933),
            .in2(N__29927),
            .in3(N__32891),
            .lcout(\this_vga_signals.g0_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_7_LC_17_19_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_7_LC_17_19_0  (
            .in0(N__29924),
            .in1(N__29918),
            .in2(N__30149),
            .in3(N__29981),
            .lcout(\this_vga_signals.if_N_10_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_7_LC_17_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_7_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_7_LC_17_19_1 .LUT_INIT=16'b1011110101000010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_7_LC_17_19_1  (
            .in0(N__31528),
            .in1(N__30565),
            .in2(N__30487),
            .in3(N__31664),
            .lcout(\this_vga_signals.g0_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_19_2 .LUT_INIT=16'b0001011100101011;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_19_2  (
            .in0(N__31666),
            .in1(N__33877),
            .in2(N__31422),
            .in3(N__30282),
            .lcout(\this_vga_signals.mult1_un61_sum_c2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_17_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_17_19_3 .LUT_INIT=16'b1101010000101011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_17_19_3  (
            .in0(N__31527),
            .in1(N__30564),
            .in2(N__30486),
            .in3(N__31663),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3 ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_N_3L3_1_LC_17_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_3L3_1_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_3L3_1_LC_17_19_4 .LUT_INIT=16'b0011001101100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_N_3L3_1_LC_17_19_4  (
            .in0(N__29900),
            .in1(N__31751),
            .in2(N__29894),
            .in3(N__30182),
            .lcout(\this_vga_signals.g0_41_N_3L3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_17_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_17_19_5 .LUT_INIT=16'b0111101100110011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_17_19_5  (
            .in0(N__33875),
            .in1(N__31526),
            .in2(N__33168),
            .in3(N__30563),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_c3_x0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_17_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_17_19_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__31037),
            .in2(N__30008),
            .in3(N__30131),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0),
            .ltout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_1_LC_17_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_1_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_41_N_4L5_1_LC_17_19_7 .LUT_INIT=16'b0001010001110010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_41_N_4L5_1_LC_17_19_7  (
            .in0(N__33876),
            .in1(N__31412),
            .in2(N__30005),
            .in3(N__31665),
            .lcout(\this_vga_signals.g0_41_N_4L5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam m31_0_x3_LC_17_20_0.C_ON=1'b0;
    defparam m31_0_x3_LC_17_20_0.SEQ_MODE=4'b0000;
    defparam m31_0_x3_LC_17_20_0.LUT_INIT=16'b0101101001011010;
    LogicCell40 m31_0_x3_LC_17_20_0 (
            .in0(N__30281),
            .in1(_gnd_net_),
            .in2(N__30413),
            .in3(_gnd_net_),
            .lcout(N_6_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_17_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_1_LC_17_20_1 .LUT_INIT=16'b0110001111011100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_1_LC_17_20_1  (
            .in0(N__30317),
            .in1(N__31754),
            .in2(N__30635),
            .in3(N__30229),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_LC_17_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_LC_17_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_LC_17_20_2  (
            .in0(N__31409),
            .in1(N__31294),
            .in2(N__29990),
            .in3(N__29987),
            .lcout(\this_vga_signals.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_17_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_0_1_LC_17_20_3 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_0_1_LC_17_20_3  (
            .in0(N__29975),
            .in1(N__30228),
            .in2(N__30038),
            .in3(N__31753),
            .lcout(),
            .ltout(\this_vga_signals.g1_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_i_o4_LC_17_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_i_o4_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_i_o4_LC_17_20_4 .LUT_INIT=16'b1000111011101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_i_o4_LC_17_20_4  (
            .in0(N__31408),
            .in1(N__31293),
            .in2(N__29969),
            .in3(N__30071),
            .lcout(\this_vga_signals.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_17_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_17_LC_17_20_5 .LUT_INIT=16'b0100000000100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_17_LC_17_20_5  (
            .in0(N__30596),
            .in1(N__30399),
            .in2(N__31421),
            .in3(N__30280),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_17_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_LC_17_20_6 .LUT_INIT=16'b0010000100001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_LC_17_20_6  (
            .in0(N__31145),
            .in1(N__33609),
            .in2(N__33182),
            .in3(N__33411),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_1_LC_17_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_1_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_1_LC_17_20_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_1_LC_17_20_7  (
            .in0(N__33931),
            .in1(_gnd_net_),
            .in2(N__30053),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.g0_0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIE8SF1_LC_17_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIE8SF1_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIE8SF1_LC_17_21_0 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIE8SF1_LC_17_21_0  (
            .in0(N__38267),
            .in1(N__34930),
            .in2(N__36566),
            .in3(N__34993),
            .lcout(M_last_q_RNIE8SF1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_17_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_17_21_1 .LUT_INIT=16'b0110011010010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_17_21_1  (
            .in0(N__31679),
            .in1(N__30509),
            .in2(N__30302),
            .in3(N__30323),
            .lcout(),
            .ltout(\this_vga_signals.N_5_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_RNIPQ17A7_2_LC_17_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_RNIPQ17A7_2_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_RNIPQ17A7_2_LC_17_21_2 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.M_vcounter_q_RNIPQ17A7_2_LC_17_21_2  (
            .in0(N__31274),
            .in1(N__31401),
            .in2(N__30050),
            .in3(N__30353),
            .lcout(\this_vga_signals.g1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_17_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_6_0_LC_17_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_6_0_LC_17_21_3  (
            .in0(N__33929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30026),
            .lcout(\this_vga_signals.g0_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_17_21_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_26_LC_17_21_4 .LUT_INIT=16'b0000100001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_26_LC_17_21_4  (
            .in0(N__33415),
            .in1(N__34069),
            .in2(N__33620),
            .in3(N__30602),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_17_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_17_21_5 .LUT_INIT=16'b0011010001000001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_17_21_5  (
            .in0(N__31130),
            .in1(N__33616),
            .in2(N__34075),
            .in3(N__33414),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2 ),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_17_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_0_LC_17_21_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_0_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30020),
            .in3(N__33928),
            .lcout(\this_vga_signals.g0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_1_LC_17_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_1_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_i_x2_1_LC_17_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_i_x2_1_LC_17_21_7  (
            .in0(N__31400),
            .in1(N__31273),
            .in2(_gnd_net_),
            .in3(N__31529),
            .lcout(\this_vga_signals.g0_i_x2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIE5RF1_LC_17_23_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIE5RF1_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIE5RF1_LC_17_23_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIE5RF1_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__36550),
            .in2(_gnd_net_),
            .in3(N__36104),
            .lcout(N_295),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_30_2.C_ON=1'b0;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_30_2.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_30_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_30_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36933),
            .lcout(GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_18_7_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_3_0_wclke_3_LC_18_7_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_spr_ram.mem_mem_3_0_wclke_3_LC_18_7_3  (
            .in0(N__32209),
            .in1(N__32116),
            .in2(N__32017),
            .in3(N__31911),
            .lcout(\this_spr_ram.mem_WE_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO4821_9_LC_18_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO4821_9_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIO4821_9_LC_18_16_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIO4821_9_LC_18_16_0  (
            .in0(N__35267),
            .in1(N__33125),
            .in2(_gnd_net_),
            .in3(N__34649),
            .lcout(\this_vga_signals.m43_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_18_16_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_18_16_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_18_16_1  (
            .in0(N__33124),
            .in1(N__33926),
            .in2(_gnd_net_),
            .in3(N__34012),
            .lcout(\this_vga_signals.vaddress_c3_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_5_LC_18_16_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_5_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_5_LC_18_16_2 .LUT_INIT=16'b1001110011000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_5_LC_18_16_2  (
            .in0(N__31522),
            .in1(N__31678),
            .in2(N__30502),
            .in3(N__30580),
            .lcout(\this_vga_signals.g0_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIKEN71_LC_18_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIKEN71_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIKEN71_LC_18_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIKEN71_LC_18_17_0  (
            .in0(N__35345),
            .in1(N__35253),
            .in2(N__34640),
            .in3(N__34729),
            .lcout(\this_vga_signals.vaddress_ac0_9_0_a0_1 ),
            .ltout(\this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNI3GK81_LC_18_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNI3GK81_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNI3GK81_LC_18_17_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNI3GK81_LC_18_17_1  (
            .in0(N__34831),
            .in1(_gnd_net_),
            .in2(N__30059),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.CO0_0_i_i ),
            .ltout(\this_vga_signals.CO0_0_i_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_0_LC_18_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_0_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_0_LC_18_17_2 .LUT_INIT=16'b1000000001001000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_0_LC_18_17_2  (
            .in0(N__32985),
            .in1(N__33121),
            .in2(N__30056),
            .in3(N__32930),
            .lcout(\this_vga_signals.N_7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_18_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_18_17_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_18_17_3  (
            .in0(N__34728),
            .in1(N__34622),
            .in2(_gnd_net_),
            .in3(N__35344),
            .lcout(),
            .ltout(\this_vga_signals.vaddress_c5_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_9_LC_18_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_9_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI3GK81_9_LC_18_17_4 .LUT_INIT=16'b1100110000111100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI3GK81_9_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__35252),
            .in2(N__30161),
            .in3(N__34830),
            .lcout(\this_vga_signals.vaddress_9 ),
            .ltout(\this_vga_signals.vaddress_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_18_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_7_LC_18_17_5 .LUT_INIT=16'b0100101100000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_7_LC_18_17_5  (
            .in0(N__34833),
            .in1(N__31064),
            .in2(N__30158),
            .in3(N__32984),
            .lcout(\this_vga_signals.g1_3_0 ),
            .ltout(\this_vga_signals.g1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_24_LC_18_17_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_24_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30155),
            .in3(N__33122),
            .lcout(\this_vga_signals.N_7_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_18_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_3_LC_18_17_7 .LUT_INIT=16'b0100101100000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_3_LC_18_17_7  (
            .in0(N__34832),
            .in1(N__31065),
            .in2(N__32943),
            .in3(N__32986),
            .lcout(\this_vga_signals.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_18_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_21_LC_18_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_21_LC_18_18_0  (
            .in0(N__31752),
            .in1(N__30283),
            .in2(_gnd_net_),
            .in3(N__31671),
            .lcout(),
            .ltout(\this_vga_signals.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_19_LC_18_18_1 .LUT_INIT=16'b1101111100000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_19_LC_18_18_1  (
            .in0(N__31407),
            .in1(N__30140),
            .in2(N__30152),
            .in3(N__30167),
            .lcout(\this_vga_signals.mult1_un61_sum_c3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_18_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_20_LC_18_18_2 .LUT_INIT=16'b0011100110011100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_20_LC_18_18_2  (
            .in0(N__31498),
            .in1(N__30403),
            .in2(N__30498),
            .in3(N__30562),
            .lcout(\this_vga_signals.N_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_18_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_18_18_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__33261),
            .in2(N__31172),
            .in3(N__31178),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_ns ),
            .ltout(\this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_18_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_18_18_4 .LUT_INIT=16'b0010000011111010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_18_18_4  (
            .in0(N__33873),
            .in1(N__33079),
            .in2(N__30134),
            .in3(N__31496),
            .lcout(\this_vga_signals.mult1_un54_sum_c3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_16_LC_18_18_5 .LUT_INIT=16'b0100000100001001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_16_LC_18_18_5  (
            .in0(N__33612),
            .in1(N__30689),
            .in2(N__33120),
            .in3(N__33407),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_18_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_18_18_6 .LUT_INIT=16'b0001101010111011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_18_18_6  (
            .in0(N__33874),
            .in1(N__31033),
            .in2(N__33149),
            .in3(N__30560),
            .lcout(\this_vga_signals.mult1_un54_sum_c2_0 ),
            .ltout(\this_vga_signals.mult1_un54_sum_c2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_18_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_40_LC_18_18_7 .LUT_INIT=16'b0000010110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_40_LC_18_18_7  (
            .in0(N__30561),
            .in1(_gnd_net_),
            .in2(N__30188),
            .in3(N__31497),
            .lcout(\this_vga_signals.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_18_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_1_LC_18_19_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_1_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__31719),
            .in2(_gnd_net_),
            .in3(N__31662),
            .lcout(),
            .ltout(\this_vga_signals.g1_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_18_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_34_LC_18_19_1 .LUT_INIT=16'b0000100000100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_34_LC_18_19_1  (
            .in0(N__31411),
            .in1(N__30393),
            .in2(N__30185),
            .in3(N__30276),
            .lcout(\this_vga_signals.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_5_LC_18_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_5_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_5_LC_18_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_5_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__31718),
            .in2(_gnd_net_),
            .in3(N__31660),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_18_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_38_LC_18_19_3 .LUT_INIT=16'b0000100000100000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_38_LC_18_19_3  (
            .in0(N__31410),
            .in1(N__30392),
            .in2(N__30176),
            .in3(N__30275),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_18_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_18_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_18_19_4  (
            .in0(N__31043),
            .in1(N__31076),
            .in2(_gnd_net_),
            .in3(N__30557),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_18_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_0_LC_18_19_5 .LUT_INIT=16'b0011111100010101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_0_LC_18_19_5  (
            .in0(N__31720),
            .in1(N__30173),
            .in2(N__30338),
            .in3(N__30227),
            .lcout(\this_vga_signals.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_5_N_2L1_LC_18_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_5_N_2L1_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_5_N_2L1_LC_18_19_6 .LUT_INIT=16'b0010101111010100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_5_N_2L1_LC_18_19_6  (
            .in0(N__31499),
            .in1(N__30559),
            .in2(N__30503),
            .in3(N__31661),
            .lcout(\this_vga_signals.g0_5_5_N_2L1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_18_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_18_19_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_18_19_7  (
            .in0(N__30558),
            .in1(N__33595),
            .in2(N__33927),
            .in3(N__31793),
            .lcout(this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_3_LC_18_20_0 .LUT_INIT=16'b0011010001000001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_3_LC_18_20_0  (
            .in0(N__31129),
            .in1(N__33614),
            .in2(N__34076),
            .in3(N__33412),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_1_LC_18_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_1_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_1_LC_18_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_1_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__31736),
            .in2(_gnd_net_),
            .in3(N__31677),
            .lcout(),
            .ltout(\this_vga_signals.g0_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_28_LC_18_20_2 .LUT_INIT=16'b0000100001000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_28_LC_18_20_2  (
            .in0(N__30279),
            .in1(N__31426),
            .in2(N__30326),
            .in3(N__30398),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_18_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_39_LC_18_20_3 .LUT_INIT=16'b0010000001000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_39_LC_18_20_3  (
            .in0(N__30397),
            .in1(N__31604),
            .in2(N__31427),
            .in3(N__30278),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_4_LC_18_20_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_4_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_4_LC_18_20_4 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_4_LC_18_20_4  (
            .in0(N__31737),
            .in1(N__31807),
            .in2(N__30311),
            .in3(N__30221),
            .lcout(\this_vga_signals.g0_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_5_LC_18_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_5_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_5_LC_18_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_5_LC_18_20_5  (
            .in0(N__30220),
            .in1(N__30293),
            .in2(N__30412),
            .in3(N__30277),
            .lcout(\this_vga_signals.g0_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_18_20_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_0_LC_18_20_6 .LUT_INIT=16'b1111001101010001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_0_LC_18_20_6  (
            .in0(N__31735),
            .in1(N__30236),
            .in2(N__31808),
            .in3(N__30219),
            .lcout(),
            .ltout(\this_vga_signals.g0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_18_20_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_4_LC_18_20_7 .LUT_INIT=16'b0110010110011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_4_LC_18_20_7  (
            .in0(N__30665),
            .in1(N__30656),
            .in2(N__30650),
            .in3(N__31676),
            .lcout(\this_vga_signals.N_5_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_1_LC_18_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_1_LC_18_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_1_LC_18_21_0 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_1_LC_18_21_0  (
            .in0(N__31524),
            .in1(N__31289),
            .in2(_gnd_net_),
            .in3(N__30582),
            .lcout(\this_vga_signals.g0_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_18_21_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_18_21_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_22_LC_18_21_1 .LUT_INIT=16'b0011010001000001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_22_LC_18_21_1  (
            .in0(N__30647),
            .in1(N__33615),
            .in2(N__34074),
            .in3(N__33416),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_18_21_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_18_21_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_LC_18_21_2 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_LC_18_21_2  (
            .in0(_gnd_net_),
            .in1(N__33930),
            .in2(N__30638),
            .in3(N__32252),
            .lcout(\this_vga_signals.g3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_18_21_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_18_21_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_33_LC_18_21_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_33_LC_18_21_3  (
            .in0(N__33105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30619),
            .lcout(\this_vga_signals.N_7_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_18_21_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_1_2_LC_18_21_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_1_2_LC_18_21_5  (
            .in0(N__31721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31675),
            .lcout(\this_vga_signals.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_18_21_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_1_LC_18_21_6 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_1_LC_18_21_6  (
            .in0(N__31525),
            .in1(N__30499),
            .in2(_gnd_net_),
            .in3(N__30583),
            .lcout(\this_vga_signals.g1_0 ),
            .ltout(\this_vga_signals.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_18_21_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_18_21_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_29_LC_18_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_29_LC_18_21_7  (
            .in0(N__30500),
            .in1(N__30428),
            .in2(N__30422),
            .in3(N__30418),
            .lcout(\this_vga_signals.g0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_7_LC_18_23_0 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_7_LC_18_23_0 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_7_LC_18_23_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_7_LC_18_23_0  (
            .in0(N__30798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30347),
            .lcout(\this_reset_cond.M_stage_qZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39369),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_9_LC_18_23_3 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_9_LC_18_23_3 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_9_LC_18_23_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \this_reset_cond.M_stage_q_9_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__30800),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(M_this_reset_cond_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39369),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_reset_cond.M_stage_q_8_LC_18_23_4 .C_ON=1'b0;
    defparam \this_reset_cond.M_stage_q_8_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \this_reset_cond.M_stage_q_8_LC_18_23_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \this_reset_cond.M_stage_q_8_LC_18_23_4  (
            .in0(N__30799),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30734),
            .lcout(\this_reset_cond.M_stage_qZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39369),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_19_7_3 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_19_7_3 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_2_0_wclke_3_LC_19_7_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \this_spr_ram.mem_mem_2_0_wclke_3_LC_19_7_3  (
            .in0(N__32217),
            .in1(N__31912),
            .in2(N__32031),
            .in3(N__32117),
            .lcout(\this_spr_ram.mem_WE_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_19_16_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_19_16_0 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_4_LC_19_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_4_LC_19_16_0  (
            .in0(N__33688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39322),
            .ce(N__34491),
            .sr(N__34428));
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_16_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_16_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_6_LC_19_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_6_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34539),
            .lcout(this_vga_signals_M_vcounter_q_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39322),
            .ce(N__34491),
            .sr(N__34428));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_16_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_16_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31572),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39322),
            .ce(N__34491),
            .sr(N__34428));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_7_LC_19_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_7_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_7_LC_19_17_0 .LUT_INIT=16'b1110111110011100;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_7_LC_19_17_0  (
            .in0(N__34837),
            .in1(N__31082),
            .in2(N__31070),
            .in3(N__32942),
            .lcout(\this_vga_signals.N_12_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_19_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_19_17_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_19_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30683),
            .in3(N__30674),
            .lcout(\this_vga_signals.vaddress_c2 ),
            .ltout(\this_vga_signals.vaddress_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_19_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_19_17_2 .LUT_INIT=16'b1010101010101001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_19_17_2  (
            .in0(N__34626),
            .in1(N__33980),
            .in2(N__30668),
            .in3(N__34730),
            .lcout(\this_vga_signals.vaddress_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_19_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_27_LC_19_17_3 .LUT_INIT=16'b0101001000100001;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_27_LC_19_17_3  (
            .in0(N__33613),
            .in1(N__31122),
            .in2(N__34017),
            .in3(N__33384),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_19_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_5_LC_19_17_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_5_LC_19_17_4  (
            .in0(N__31103),
            .in1(_gnd_net_),
            .in2(N__31097),
            .in3(N__33939),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0_6_LC_19_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0_6_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0_6_LC_19_17_5 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0_6_LC_19_17_5  (
            .in0(N__35184),
            .in1(N__35313),
            .in2(N__32861),
            .in3(N__32882),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_19_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_19_17_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_19_17_6  (
            .in0(N__35312),
            .in1(N__32856),
            .in2(_gnd_net_),
            .in3(N__35183),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_7_LC_19_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_7_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNI65531_0_7_LC_19_17_7 .LUT_INIT=16'b0011001100110110;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNI65531_0_7_LC_19_17_7  (
            .in0(N__34731),
            .in1(N__34627),
            .in2(N__34016),
            .in3(N__34836),
            .lcout(\this_vga_signals.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_19_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_19_18_0 .LUT_INIT=16'b0010010011011011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_19_18_0  (
            .in0(N__33479),
            .in1(N__33440),
            .in2(N__33254),
            .in3(N__31781),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_19_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_19_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g1_5_LC_19_18_1 .LUT_INIT=16'b0010001010010010;
    LogicCell40 \this_vga_signals.un5_vaddress_g1_5_LC_19_18_1  (
            .in0(N__32983),
            .in1(N__32929),
            .in2(N__31069),
            .in3(N__34835),
            .lcout(\this_vga_signals.g1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_19_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_19_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_19_18_2 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_19_18_2  (
            .in0(N__33478),
            .in1(N__33442),
            .in2(N__33253),
            .in3(N__31782),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc3_1_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_19_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_19_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_19_18_3 .LUT_INIT=16'b0011110001011010;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_19_18_3  (
            .in0(N__31783),
            .in1(N__33238),
            .in2(N__31598),
            .in3(N__33295),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_19_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_19_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_19_18_4 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_19_18_4  (
            .in0(N__33237),
            .in1(N__33474),
            .in2(_gnd_net_),
            .in3(N__33441),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34_6_LC_19_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34_6_LC_19_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34_6_LC_19_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34_6_LC_19_18_5  (
            .in0(N__31451),
            .in1(N__31445),
            .in2(_gnd_net_),
            .in3(N__34834),
            .lcout(),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1_6_LC_19_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1_6_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1_6_LC_19_18_6 .LUT_INIT=16'b1001011001100110;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1_6_LC_19_18_6  (
            .in0(N__33532),
            .in1(N__33473),
            .in2(N__31439),
            .in3(N__32831),
            .lcout(\this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6 ),
            .ltout(\this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x0_LC_19_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x0_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x0_LC_19_18_7 .LUT_INIT=16'b1001100101101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x0_LC_19_18_7  (
            .in0(N__31594),
            .in1(N__33901),
            .in2(N__31436),
            .in3(N__33294),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_42_LC_19_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_42_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_42_LC_19_19_0 .LUT_INIT=16'b0110010110100110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_42_LC_19_19_0  (
            .in0(N__31433),
            .in1(N__31399),
            .in2(N__31295),
            .in3(N__31193),
            .lcout(\this_vga_signals.N_5786_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_19_19_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_19_19_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_19_19_1 .LUT_INIT=16'b0000000010010110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_19_19_1  (
            .in0(N__33475),
            .in1(N__33358),
            .in2(N__33573),
            .in3(N__33292),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_x0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_19_19_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_19_19_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_19_19_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_19_19_2  (
            .in0(N__33293),
            .in1(N__33356),
            .in2(N__33572),
            .in3(N__33476),
            .lcout(\this_vga_signals.mult1_un47_sum_axbxc3_x1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_0_7_LC_19_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_0_7_LC_19_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_0_7_LC_19_19_3 .LUT_INIT=16'b0111011110011001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_0_7_LC_19_19_3  (
            .in0(N__31163),
            .in1(N__33001),
            .in2(_gnd_net_),
            .in3(N__32944),
            .lcout(\this_vga_signals.N_12_0 ),
            .ltout(\this_vga_signals.N_12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_0_LC_19_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_0_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_0_LC_19_19_4 .LUT_INIT=16'b0100000000100101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_0_LC_19_19_4  (
            .in0(N__33536),
            .in1(N__33357),
            .in2(N__31133),
            .in3(N__33083),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_1_LC_19_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_1_LC_19_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_1_LC_19_19_5 .LUT_INIT=16'b0111000110001110;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_1_LC_19_19_5  (
            .in0(N__33477),
            .in1(N__33443),
            .in2(N__33266),
            .in3(N__33359),
            .lcout(\this_vga_signals.mult1_un61_sum_axb1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_19_7 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_5_LC_19_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_5_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31573),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39345),
            .ce(N__34509),
            .sr(N__34430));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x1_LC_19_20_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x1_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x1_LC_19_20_0 .LUT_INIT=16'b0101101001101001;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x1_LC_19_20_0  (
            .in0(N__31593),
            .in1(N__31787),
            .in2(N__33943),
            .in3(N__33296),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_ns_LC_19_20_1 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_ns_LC_19_20_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_ns_LC_19_20_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_ns_LC_19_20_1  (
            .in0(N__33265),
            .in1(_gnd_net_),
            .in2(N__31766),
            .in3(N__31763),
            .lcout(\this_vga_signals.mult1_un54_sum_axbxc1_ns ),
            .ltout(\this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_19_20_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_19_20_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_2_2_LC_19_20_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_2_2_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31682),
            .in3(N__31667),
            .lcout(\this_vga_signals.g0_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_0_LC_19_20_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_0_LC_19_20_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_0_LC_19_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_0_LC_19_20_3  (
            .in0(_gnd_net_),
            .in1(N__33640),
            .in2(_gnd_net_),
            .in3(N__33659),
            .lcout(\this_vga_signals.mult1_un54_sum_axb1_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_20_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_20_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31577),
            .lcout(\this_vga_signals.M_vcounter_q_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39354),
            .ce(N__34510),
            .sr(N__34432));
    defparam \this_start_data_delay.M_last_q_RNI1KH61_LC_19_21_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI1KH61_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI1KH61_LC_19_21_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI1KH61_LC_19_21_0  (
            .in0(N__31550),
            .in1(N__35539),
            .in2(N__33701),
            .in3(N__36616),
            .lcout(\this_start_data_delay.N_380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_19_21_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_19_21_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_start_data_delay.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_19_21_2  (
            .in0(N__34327),
            .in1(N__34350),
            .in2(N__33776),
            .in3(N__34367),
            .lcout(),
            .ltout(M_this_state_d_0_sqmuxa_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_substate_q_LC_19_21_3.C_ON=1'b0;
    defparam M_this_substate_q_LC_19_21_3.SEQ_MODE=4'b1000;
    defparam M_this_substate_q_LC_19_21_3.LUT_INIT=16'b1110001010101010;
    LogicCell40 M_this_substate_q_LC_19_21_3 (
            .in0(N__34368),
            .in1(N__38007),
            .in2(N__32300),
            .in3(N__35921),
            .lcout(M_this_substate_qZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39362),
            .ce(),
            .sr(N__36812));
    defparam \this_start_data_delay.M_last_q_RNIO2A13_0_LC_19_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIO2A13_0_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIO2A13_0_LC_19_21_5 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \this_start_data_delay.M_last_q_RNIO2A13_0_LC_19_21_5  (
            .in0(N__36617),
            .in1(N__38334),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\this_start_data_delay.N_233_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIHUID5_LC_19_21_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIHUID5_LC_19_21_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIHUID5_LC_19_21_6 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \this_start_data_delay.M_last_q_RNIHUID5_LC_19_21_6  (
            .in0(N__35909),
            .in1(N__37045),
            .in2(N__32297),
            .in3(N__36935),
            .lcout(N_164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_19_22_3 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_19_22_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_23_LC_19_22_3 .LUT_INIT=16'b0001010000000110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_23_LC_19_22_3  (
            .in0(N__33594),
            .in1(N__32264),
            .in2(N__33131),
            .in3(N__33413),
            .lcout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICPQ11_LC_19_23_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICPQ11_LC_19_23_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICPQ11_LC_19_23_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNICPQ11_LC_19_23_3  (
            .in0(_gnd_net_),
            .in1(N__36565),
            .in2(_gnd_net_),
            .in3(N__36134),
            .lcout(N_93),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_1_3_LC_19_24_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_1_3_LC_19_24_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_1_3_LC_19_24_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_1_3_LC_19_24_0  (
            .in0(N__35426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35469),
            .lcout(\this_start_data_delay.N_467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_20_11_4 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_4_0_wclke_3_LC_20_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \this_spr_ram.mem_mem_4_0_wclke_3_LC_20_11_4  (
            .in0(N__32205),
            .in1(N__32103),
            .in2(N__32016),
            .in3(N__31918),
            .lcout(\this_spr_ram.mem_WE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_20_13_0 .C_ON=1'b0;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_20_13_0 .SEQ_MODE=4'b0000;
    defparam \this_spr_ram.mem_mem_5_0_wclke_3_LC_20_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \this_spr_ram.mem_mem_5_0_wclke_3_LC_20_13_0  (
            .in0(N__32177),
            .in1(N__32081),
            .in2(N__31996),
            .in3(N__31913),
            .lcout(\this_spr_ram.mem_WE_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIPTJA2_LC_20_15_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIPTJA2_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIPTJA2_LC_20_15_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIPTJA2_LC_20_15_4  (
            .in0(N__37891),
            .in1(N__35131),
            .in2(N__38737),
            .in3(N__38278),
            .lcout(M_this_spr_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_20_16_1 .C_ON=1'b0;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_20_16_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_20_16_1  (
            .in0(N__32735),
            .in1(N__32723),
            .in2(_gnd_net_),
            .in3(N__32693),
            .lcout(M_this_ppu_spr_addr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_0_12_LC_20_16_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_0_12_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_0_12_LC_20_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_0_12_LC_20_16_5  (
            .in0(_gnd_net_),
            .in1(N__38348),
            .in2(_gnd_net_),
            .in3(N__35712),
            .lcout(\this_start_data_delay.N_284_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNILPJA2_LC_20_16_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNILPJA2_LC_20_16_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNILPJA2_LC_20_16_7 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNILPJA2_LC_20_16_7  (
            .in0(N__37766),
            .in1(N__35130),
            .in2(N__38896),
            .in3(N__38281),
            .lcout(M_this_spr_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_6_LC_20_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_6_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_6_LC_20_17_0 .LUT_INIT=16'b1111011100001111;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_6_LC_20_17_0  (
            .in0(N__35180),
            .in1(N__32879),
            .in2(N__32860),
            .in3(N__35306),
            .lcout(\this_vga_signals.m47_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_20_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_6_LC_20_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_6_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34546),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39337),
            .ce(N__34498),
            .sr(N__34429));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34564),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39337),
            .ce(N__34498),
            .sr(N__34429));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34771),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39337),
            .ce(N__34498),
            .sr(N__34429));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34672),
            .lcout(\this_vga_signals.M_vcounter_q_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39337),
            .ce(N__34498),
            .sr(N__34429));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_1_LC_20_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_1_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_1_LC_20_17_5 .LUT_INIT=16'b0100111100001100;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_1_LC_20_17_5  (
            .in0(N__32880),
            .in1(N__32854),
            .in2(N__35189),
            .in3(N__35314),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_20_17_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_20_17_6 .LUT_INIT=16'b1010011111110101;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_20_17_6  (
            .in0(N__35230),
            .in1(N__34828),
            .in2(N__33272),
            .in3(N__35307),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_17_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_17_7 .LUT_INIT=16'b1011000011010000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_17_7  (
            .in0(N__34829),
            .in1(N__34628),
            .in2(N__33269),
            .in3(N__35150),
            .lcout(\this_vga_signals.mult1_un40_sum_c3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_20_18_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_30_LC_20_18_0 .LUT_INIT=16'b0000010000011010;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_30_LC_20_18_0  (
            .in0(N__33194),
            .in1(N__33380),
            .in2(N__33582),
            .in3(N__33078),
            .lcout(),
            .ltout(\this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9FPA_4_LC_20_18_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9FPA_4_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIE9FPA_4_LC_20_18_1 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIE9FPA_4_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(N__33903),
            .in2(N__33212),
            .in3(N__33008),
            .lcout(\this_vga_signals.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_20_18_2 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_35_LC_20_18_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_35_LC_20_18_2  (
            .in0(N__33193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33077),
            .lcout(),
            .ltout(\this_vga_signals.N_7_1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLNC5_6_LC_20_18_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLNC5_6_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_esr_RNIOLNC5_6_LC_20_18_3 .LUT_INIT=16'b0010011000001001;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_RNIOLNC5_6_LC_20_18_3  (
            .in0(N__34019),
            .in1(N__33546),
            .in2(N__33011),
            .in3(N__33370),
            .lcout(\this_vga_signals.G_5_i_o2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_20_18_4 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_32_LC_20_18_4 .LUT_INIT=16'b1010001000101000;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_32_LC_20_18_4  (
            .in0(N__33782),
            .in1(N__32996),
            .in2(N__34784),
            .in3(N__32948),
            .lcout(\this_vga_signals.N_19_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_1_6_LC_20_18_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_1_6_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_1_6_LC_20_18_5 .LUT_INIT=16'b0011000001000101;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_1_6_LC_20_18_5  (
            .in0(N__32881),
            .in1(N__32855),
            .in2(N__35315),
            .in3(N__35181),
            .lcout(),
            .ltout(\this_vga_signals.m47_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIDJ05_7_LC_20_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIDJ05_7_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_fast_esr_RNIDJ05_7_LC_20_18_6 .LUT_INIT=16'b0100110010001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_fast_esr_RNIDJ05_7_LC_20_18_6  (
            .in0(N__35182),
            .in1(N__32830),
            .in2(N__34079),
            .in3(N__34827),
            .lcout(\this_vga_signals.SUM_2 ),
            .ltout(\this_vga_signals.SUM_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a7_1_3_LC_20_18_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a7_1_3_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_a7_1_3_LC_20_18_7 .LUT_INIT=16'b0100000000000100;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_a7_1_3_LC_20_18_7  (
            .in0(N__34018),
            .in1(N__33902),
            .in2(N__33785),
            .in3(N__33545),
            .lcout(\this_vga_signals.g0_0_i_a7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_LC_20_19_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_LC_20_19_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \this_vga_signals.M_this_state_d28_0_a2_0_LC_20_19_0  (
            .in0(N__33719),
            .in1(N__33764),
            .in2(N__33746),
            .in3(N__35540),
            .lcout(N_88),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1_6_LC_20_19_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1_6_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1_6_LC_20_19_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1_6_LC_20_19_1  (
            .in0(N__33763),
            .in1(N__33742),
            .in2(_gnd_net_),
            .in3(N__33718),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_19_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(N__33635),
            .in2(_gnd_net_),
            .in3(N__33657),
            .lcout(\this_vga_signals.vaddress_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_20_19_4 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_20_19_4 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_20_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_20_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33689),
            .lcout(\this_vga_signals.M_vcounter_q_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39355),
            .ce(N__34511),
            .sr(N__34433));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_20_19_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_20_19_5 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_20_19_5  (
            .in0(N__35342),
            .in1(N__33636),
            .in2(_gnd_net_),
            .in3(N__33656),
            .lcout(\this_vga_signals.vaddress_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI88ES_LC_20_19_6 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI88ES_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI88ES_LC_20_19_6 .LUT_INIT=16'b1100110010010011;
    LogicCell40 \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI88ES_LC_20_19_6  (
            .in0(N__33658),
            .in1(N__34733),
            .in2(N__33641),
            .in3(N__35343),
            .lcout(\this_vga_signals.vaddress_7 ),
            .ltout(\this_vga_signals.vaddress_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_m2_0_LC_20_19_7 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_m2_0_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_m2_0_LC_20_19_7 .LUT_INIT=16'b0000011001100000;
    LogicCell40 \this_vga_signals.un5_vaddress_if_m2_0_LC_20_19_7  (
            .in0(N__33472),
            .in1(N__33439),
            .in2(N__33419),
            .in3(N__33355),
            .lcout(\this_vga_signals.if_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIK6R81_0_LC_20_20_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_0_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIK6R81_0_LC_20_20_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIK6R81_0_LC_20_20_0  (
            .in0(N__35607),
            .in1(N__38229),
            .in2(_gnd_net_),
            .in3(N__36562),
            .lcout(\this_start_data_delay.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIGR6G1_LC_20_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIGR6G1_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIGR6G1_LC_20_20_1 .LUT_INIT=16'b0011000000010000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIGR6G1_LC_20_20_1  (
            .in0(N__36563),
            .in1(N__36953),
            .in2(N__36035),
            .in3(N__37997),
            .lcout(),
            .ltout(\this_start_data_delay.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_1_LC_20_20_2.C_ON=1'b0;
    defparam M_this_state_q_1_LC_20_20_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_1_LC_20_20_2.LUT_INIT=16'b1111000111110000;
    LogicCell40 M_this_state_q_1_LC_20_20_2 (
            .in0(N__35417),
            .in1(N__35476),
            .in2(N__34100),
            .in3(N__35363),
            .lcout(M_this_state_qZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39363),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIH1242_LC_20_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIH1242_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIH1242_LC_20_20_6 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIH1242_LC_20_20_6  (
            .in0(N__36952),
            .in1(N__36564),
            .in2(N__35713),
            .in3(N__36632),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_12_LC_20_20_7.C_ON=1'b0;
    defparam M_this_state_q_12_LC_20_20_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_12_LC_20_20_7.LUT_INIT=16'b1111000011100000;
    LogicCell40 M_this_state_q_12_LC_20_20_7 (
            .in0(N__34097),
            .in1(N__36166),
            .in2(N__34088),
            .in3(N__34903),
            .lcout(M_this_state_qZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39363),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_6_LC_20_21_0.C_ON=1'b0;
    defparam M_this_state_q_6_LC_20_21_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_6_LC_20_21_0.LUT_INIT=16'b1110110010100000;
    LogicCell40 M_this_state_q_6_LC_20_21_0 (
            .in0(N__34301),
            .in1(N__35963),
            .in2(N__34379),
            .in3(N__36165),
            .lcout(M_this_state_qZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39370),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINO621_LC_20_21_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINO621_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINO621_LC_20_21_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.M_last_q_RNINO621_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(N__36568),
            .in2(_gnd_net_),
            .in3(N__36937),
            .lcout(\this_start_data_delay.N_23_1_0 ),
            .ltout(\this_start_data_delay.N_23_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIMS691_LC_20_21_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIMS691_LC_20_21_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIMS691_LC_20_21_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIMS691_LC_20_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34085),
            .in3(N__36086),
            .lcout(),
            .ltout(\this_start_data_delay.N_339_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_3_LC_20_21_3.C_ON=1'b0;
    defparam M_this_state_q_3_LC_20_21_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_3_LC_20_21_3.LUT_INIT=16'b1111100011110000;
    LogicCell40 M_this_state_q_3_LC_20_21_3 (
            .in0(N__34352),
            .in1(N__34370),
            .in2(N__34082),
            .in3(N__35366),
            .lcout(M_this_state_qZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39370),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1_6_LC_20_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1_6_LC_20_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1_6_LC_20_21_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1_6_LC_20_21_4  (
            .in0(N__36938),
            .in1(N__34326),
            .in2(N__35507),
            .in3(N__37979),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIGTHM1_LC_20_21_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIGTHM1_LC_20_21_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIGTHM1_LC_20_21_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIGTHM1_LC_20_21_5  (
            .in0(N__37978),
            .in1(N__34299),
            .in2(N__34328),
            .in3(N__36939),
            .lcout(\this_start_data_delay.N_386 ),
            .ltout(\this_start_data_delay.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_2_LC_20_21_6.C_ON=1'b0;
    defparam M_this_state_q_2_LC_20_21_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_2_LC_20_21_6.LUT_INIT=16'b1111111101000000;
    LogicCell40 M_this_state_q_2_LC_20_21_6 (
            .in0(N__34369),
            .in1(N__34351),
            .in2(N__34331),
            .in3(N__34289),
            .lcout(M_this_state_qZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39370),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_21_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_21_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_21_7 .LUT_INIT=16'b0100010011000100;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_21_7  (
            .in0(N__34325),
            .in1(N__34300),
            .in2(N__35424),
            .in3(N__35459),
            .lcout(N_465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_22_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNILR691_LC_20_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNILR691_LC_20_22_2  (
            .in0(_gnd_net_),
            .in1(N__35961),
            .in2(_gnd_net_),
            .in3(N__36055),
            .lcout(\this_start_data_delay.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNINRJA2_LC_21_15_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNINRJA2_LC_21_15_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNINRJA2_LC_21_15_3 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNINRJA2_LC_21_15_3  (
            .in0(N__37651),
            .in1(N__35135),
            .in2(N__37331),
            .in3(N__38279),
            .lcout(M_this_spr_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_0_LC_21_16_1 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_0_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_0_LC_21_16_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_0_a2_0_LC_21_16_1  (
            .in0(N__35726),
            .in1(N__36593),
            .in2(N__34916),
            .in3(N__35660),
            .lcout(),
            .ltout(dma_axb0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dma_c4_LC_21_16_2.C_ON=1'b0;
    defparam dma_c4_LC_21_16_2.SEQ_MODE=4'b0000;
    defparam dma_c4_LC_21_16_2.LUT_INIT=16'b1111111000000000;
    LogicCell40 dma_c4_LC_21_16_2 (
            .in0(N__34850),
            .in1(N__34940),
            .in2(N__34181),
            .in3(N__34106),
            .lcout(dma_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_LC_21_16_5 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_LC_21_16_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_LC_21_16_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_3_LC_21_16_5  (
            .in0(N__35611),
            .in1(N__38280),
            .in2(_gnd_net_),
            .in3(N__35144),
            .lcout(dma_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_g0_0_i_o2_0_LC_21_17_0 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_o2_0_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_g0_0_i_o2_0_LC_21_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \this_vga_signals.un5_vaddress_g0_0_i_o2_0_LC_21_17_0  (
            .in0(N__35239),
            .in1(N__34716),
            .in2(N__34632),
            .in3(N__34841),
            .lcout(\this_vga_signals.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_17_1 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_17_1 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_7_LC_21_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_7_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34775),
            .lcout(this_vga_signals_M_vcounter_q_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39346),
            .ce(N__34508),
            .sr(N__34431));
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_17_2 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_17_2 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_8_LC_21_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_8_LC_21_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34676),
            .lcout(this_vga_signals_M_vcounter_q_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39346),
            .ce(N__34508),
            .sr(N__34431));
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_17_3 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_17_3 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_esr_9_LC_21_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_esr_9_LC_21_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34568),
            .lcout(\this_vga_signals.M_vcounter_qZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39346),
            .ce(N__34508),
            .sr(N__34431));
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_21_17_5 .C_ON=1'b0;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_21_17_5 .SEQ_MODE=4'b1000;
    defparam \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_21_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_21_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34547),
            .lcout(\this_vga_signals.M_vcounter_q_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39346),
            .ce(N__34508),
            .sr(N__34431));
    defparam M_this_state_q_13_LC_21_18_0.C_ON=1'b0;
    defparam M_this_state_q_13_LC_21_18_0.SEQ_MODE=4'b1000;
    defparam M_this_state_q_13_LC_21_18_0.LUT_INIT=16'b1010100010001000;
    LogicCell40 M_this_state_q_13_LC_21_18_0 (
            .in0(N__35972),
            .in1(N__34892),
            .in2(N__36992),
            .in3(N__35714),
            .lcout(M_this_state_qZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39356),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_11_LC_21_18_2.C_ON=1'b0;
    defparam M_this_state_q_11_LC_21_18_2.SEQ_MODE=4'b1000;
    defparam M_this_state_q_11_LC_21_18_2.LUT_INIT=16'b1010101010000000;
    LogicCell40 M_this_state_q_11_LC_21_18_2 (
            .in0(N__35971),
            .in1(N__36421),
            .in2(N__36991),
            .in3(N__34984),
            .lcout(M_this_state_qZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39356),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_6__m6_i_a4_0_a2_2_LC_21_18_4.C_ON=1'b0;
    defparam led_1_7_6__m6_i_a4_0_a2_2_LC_21_18_4.SEQ_MODE=4'b0000;
    defparam led_1_7_6__m6_i_a4_0_a2_2_LC_21_18_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 led_1_7_6__m6_i_a4_0_a2_2_LC_21_18_4 (
            .in0(N__35628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38285),
            .lcout(),
            .ltout(N_422_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_6__N_458_i_LC_21_18_5.C_ON=1'b0;
    defparam led_1_7_6__N_458_i_LC_21_18_5.SEQ_MODE=4'b0000;
    defparam led_1_7_6__N_458_i_LC_21_18_5.LUT_INIT=16'b1110111111111111;
    LogicCell40 led_1_7_6__N_458_i_LC_21_18_5 (
            .in0(N__34893),
            .in1(N__34985),
            .in2(N__34403),
            .in3(N__37939),
            .lcout(N_458_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_21_18_6 .C_ON=1'b0;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_21_18_6 .LUT_INIT=16'b0001010101010111;
    LogicCell40 \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_21_18_6  (
            .in0(N__35336),
            .in1(N__35311),
            .in2(N__35251),
            .in3(N__35185),
            .lcout(\this_vga_signals.mult1_un40_sum_ac0_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_10_LC_21_19_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_10_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_10_LC_21_19_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_10_LC_21_19_0  (
            .in0(N__34974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36130),
            .lcout(\this_start_data_delay.N_242_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_1_3_LC_21_19_3 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_1_3_LC_21_19_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_1_3_LC_21_19_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_1_3_LC_21_19_3  (
            .in0(N__35695),
            .in1(N__34973),
            .in2(N__34894),
            .in3(N__36413),
            .lcout(\this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_4_LC_21_19_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_4_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_4_LC_21_19_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_4_LC_21_19_4  (
            .in0(N__35480),
            .in1(N__35425),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.N_387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIJNJA2_LC_21_19_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIJNJA2_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIJNJA2_LC_21_19_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIJNJA2_LC_21_19_5  (
            .in0(N__38116),
            .in1(N__35120),
            .in2(N__37521),
            .in3(N__38284),
            .lcout(M_this_spr_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_o2_1_LC_21_20_0 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_o2_1_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_o2_1_LC_21_20_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_0_o2_1_LC_21_20_0  (
            .in0(_gnd_net_),
            .in1(N__36414),
            .in2(_gnd_net_),
            .in3(N__35652),
            .lcout(\this_start_data_delay.N_245_0 ),
            .ltout(\this_start_data_delay.N_245_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_1_LC_21_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_1_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_1_LC_21_20_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_0_a2_1_LC_21_20_1  (
            .in0(N__36161),
            .in1(N__34986),
            .in2(N__34943),
            .in3(N__35983),
            .lcout(un20_i_a4_0_a2_0_a2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_2_LC_21_20_2 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_2_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_2_LC_21_20_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_2_LC_21_20_2  (
            .in0(N__35710),
            .in1(N__36097),
            .in2(N__34907),
            .in3(N__35653),
            .lcout(un20_i_a4_0_a2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNICVMT3_LC_21_20_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNICVMT3_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNICVMT3_LC_21_20_3 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \this_start_data_delay.M_last_q_RNICVMT3_LC_21_20_3  (
            .in0(N__35654),
            .in1(N__36631),
            .in2(N__38141),
            .in3(N__36954),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_7_LC_21_20_4.C_ON=1'b0;
    defparam M_this_state_q_7_LC_21_20_4.SEQ_MODE=4'b1000;
    defparam M_this_state_q_7_LC_21_20_4.LUT_INIT=16'b1111000011100000;
    LogicCell40 M_this_state_q_7_LC_21_20_4 (
            .in0(N__35805),
            .in1(N__38228),
            .in2(N__35729),
            .in3(N__35655),
            .lcout(M_this_state_qZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39371),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_2_0_LC_21_20_5 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_2_0_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_0_a2_2_0_LC_21_20_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_0_a2_2_0_LC_21_20_5  (
            .in0(N__38227),
            .in1(N__36007),
            .in2(_gnd_net_),
            .in3(N__36085),
            .lcout(\this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o4_0_LC_21_20_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o4_0_LC_21_20_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_data_count_qlde_i_o4_0_LC_21_20_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \this_start_data_delay.M_this_data_count_qlde_i_o4_0_LC_21_20_6  (
            .in0(N__35711),
            .in1(_gnd_net_),
            .in2(N__35669),
            .in3(_gnd_net_),
            .lcout(\this_start_data_delay.N_246_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_8_LC_21_20_7.C_ON=1'b0;
    defparam M_this_state_q_8_LC_21_20_7.SEQ_MODE=4'b1000;
    defparam M_this_state_q_8_LC_21_20_7.LUT_INIT=16'b1100110010000000;
    LogicCell40 M_this_state_q_8_LC_21_20_7 (
            .in0(N__35656),
            .in1(N__35965),
            .in2(N__36984),
            .in3(N__35620),
            .lcout(M_this_state_qZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39371),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_1_LC_21_21_0 .C_ON=1'b0;
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_1_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \this_vga_signals.M_this_state_d28_0_a2_0_1_LC_21_21_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \this_vga_signals.M_this_state_d28_0_a2_0_1_LC_21_21_0  (
            .in0(N__35573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35558),
            .lcout(this_vga_signals_M_this_state_d28_0_a2_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_RNIKV6G1_2_LC_21_21_1.C_ON=1'b0;
    defparam M_this_state_q_RNIKV6G1_2_LC_21_21_1.SEQ_MODE=4'b0000;
    defparam M_this_state_q_RNIKV6G1_2_LC_21_21_1.LUT_INIT=16'b1010101011101010;
    LogicCell40 M_this_state_q_RNIKV6G1_2_LC_21_21_1 (
            .in0(N__36936),
            .in1(N__36084),
            .in2(N__36572),
            .in3(N__36054),
            .lcout(N_1264_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_4_LC_21_21_3.C_ON=1'b0;
    defparam M_this_state_q_4_LC_21_21_3.SEQ_MODE=4'b1000;
    defparam M_this_state_q_4_LC_21_21_3.LUT_INIT=16'b1110101011000000;
    LogicCell40 M_this_state_q_4_LC_21_21_3 (
            .in0(N__38160),
            .in1(N__35365),
            .in2(N__35503),
            .in3(N__35964),
            .lcout(M_this_state_qZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39377),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_21_21_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_21_21_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIOU691_LC_21_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIOU691_LC_21_21_4  (
            .in0(_gnd_net_),
            .in1(N__35962),
            .in2(_gnd_net_),
            .in3(N__36126),
            .lcout(),
            .ltout(\this_start_data_delay.N_337_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_5_LC_21_21_5.C_ON=1'b0;
    defparam M_this_state_q_5_LC_21_21_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_5_LC_21_21_5.LUT_INIT=16'b1111100011110000;
    LogicCell40 M_this_state_q_5_LC_21_21_5 (
            .in0(N__35460),
            .in1(N__35413),
            .in2(N__35369),
            .in3(N__35364),
            .lcout(M_this_state_qZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39377),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_ext_address_d_0_sqmuxa_1_0_a4_0_o2_i_o4_LC_21_21_6 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_ext_address_d_0_sqmuxa_1_0_a4_0_o2_i_o4_LC_21_21_6 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_ext_address_d_0_sqmuxa_1_0_a4_0_o2_i_o4_LC_21_21_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \this_start_data_delay.M_this_ext_address_d_0_sqmuxa_1_0_a4_0_o2_i_o4_LC_21_21_6  (
            .in0(N__36160),
            .in1(N__38159),
            .in2(_gnd_net_),
            .in3(N__36125),
            .lcout(\this_start_data_delay.N_239_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_0_a4_1_LC_21_21_7 .C_ON=1'b0;
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_0_a4_1_LC_21_21_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.un20_i_a4_0_a2_3_0_a4_1_LC_21_21_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \this_start_data_delay.un20_i_a4_0_a2_3_0_a4_1_LC_21_21_7  (
            .in0(_gnd_net_),
            .in1(N__36083),
            .in2(_gnd_net_),
            .in3(N__36053),
            .lcout(\this_start_data_delay.N_420_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_LC_21_22_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_LC_21_22_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_LC_21_22_4  (
            .in0(_gnd_net_),
            .in1(N__36020),
            .in2(_gnd_net_),
            .in3(N__35984),
            .lcout(N_466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIVPN44_LC_21_22_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIVPN44_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIVPN44_LC_21_22_5 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIVPN44_LC_21_22_5  (
            .in0(N__38344),
            .in1(N__35904),
            .in2(N__37996),
            .in3(N__35960),
            .lcout(),
            .ltout(\this_start_data_delay.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_0_LC_21_22_6.C_ON=1'b0;
    defparam M_this_state_q_0_LC_21_22_6.SEQ_MODE=4'b1000;
    defparam M_this_state_q_0_LC_21_22_6.LUT_INIT=16'b0000010100001101;
    LogicCell40 M_this_state_q_0_LC_21_22_6 (
            .in0(N__35885),
            .in1(N__37983),
            .in2(N__35924),
            .in3(N__35920),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39385),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_0_LC_21_22_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_0_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_0_LC_21_22_7 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_0_LC_21_22_7  (
            .in0(N__38345),
            .in1(N__35905),
            .in2(N__37938),
            .in3(N__36950),
            .lcout(\this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_ext_address_q_0_LC_21_24_0.C_ON=1'b1;
    defparam M_this_ext_address_q_0_LC_21_24_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_0_LC_21_24_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_0_LC_21_24_0 (
            .in0(N__37090),
            .in1(N__35851),
            .in2(N__35879),
            .in3(N__35878),
            .lcout(M_this_ext_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_21_24_0_),
            .carryout(un1_M_this_ext_address_q_cry_0),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_1_LC_21_24_1.C_ON=1'b1;
    defparam M_this_ext_address_q_1_LC_21_24_1.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_1_LC_21_24_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_1_LC_21_24_1 (
            .in0(N__37094),
            .in1(N__35827),
            .in2(_gnd_net_),
            .in3(N__35816),
            .lcout(M_this_ext_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_0),
            .carryout(un1_M_this_ext_address_q_cry_1),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_2_LC_21_24_2.C_ON=1'b1;
    defparam M_this_ext_address_q_2_LC_21_24_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_2_LC_21_24_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_2_LC_21_24_2 (
            .in0(N__37091),
            .in1(N__36382),
            .in2(_gnd_net_),
            .in3(N__36371),
            .lcout(M_this_ext_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_1),
            .carryout(un1_M_this_ext_address_q_cry_2),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_3_LC_21_24_3.C_ON=1'b1;
    defparam M_this_ext_address_q_3_LC_21_24_3.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_3_LC_21_24_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_3_LC_21_24_3 (
            .in0(N__37095),
            .in1(N__36355),
            .in2(_gnd_net_),
            .in3(N__36344),
            .lcout(M_this_ext_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_2),
            .carryout(un1_M_this_ext_address_q_cry_3),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_4_LC_21_24_4.C_ON=1'b1;
    defparam M_this_ext_address_q_4_LC_21_24_4.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_4_LC_21_24_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_4_LC_21_24_4 (
            .in0(N__37092),
            .in1(N__36328),
            .in2(_gnd_net_),
            .in3(N__36317),
            .lcout(M_this_ext_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_3),
            .carryout(un1_M_this_ext_address_q_cry_4),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_5_LC_21_24_5.C_ON=1'b1;
    defparam M_this_ext_address_q_5_LC_21_24_5.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_5_LC_21_24_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_5_LC_21_24_5 (
            .in0(N__37096),
            .in1(N__36301),
            .in2(_gnd_net_),
            .in3(N__36290),
            .lcout(M_this_ext_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_4),
            .carryout(un1_M_this_ext_address_q_cry_5),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_6_LC_21_24_6.C_ON=1'b1;
    defparam M_this_ext_address_q_6_LC_21_24_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_6_LC_21_24_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_6_LC_21_24_6 (
            .in0(N__37093),
            .in1(N__36271),
            .in2(_gnd_net_),
            .in3(N__36260),
            .lcout(M_this_ext_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_5),
            .carryout(un1_M_this_ext_address_q_cry_6),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_7_LC_21_24_7.C_ON=1'b1;
    defparam M_this_ext_address_q_7_LC_21_24_7.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_7_LC_21_24_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_ext_address_q_7_LC_21_24_7 (
            .in0(N__37097),
            .in1(N__36241),
            .in2(_gnd_net_),
            .in3(N__36230),
            .lcout(M_this_ext_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_6),
            .carryout(un1_M_this_ext_address_q_cry_7),
            .clk(N__39397),
            .ce(),
            .sr(N__36815));
    defparam M_this_ext_address_q_8_LC_21_25_0.C_ON=1'b1;
    defparam M_this_ext_address_q_8_LC_21_25_0.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_8_LC_21_25_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_8_LC_21_25_0 (
            .in0(N__38117),
            .in1(N__37082),
            .in2(N__36217),
            .in3(N__36200),
            .lcout(M_this_ext_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_21_25_0_),
            .carryout(un1_M_this_ext_address_q_cry_8),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_9_LC_21_25_1.C_ON=1'b1;
    defparam M_this_ext_address_q_9_LC_21_25_1.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_9_LC_21_25_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_9_LC_21_25_1 (
            .in0(N__37751),
            .in1(N__37086),
            .in2(N__36190),
            .in3(N__36173),
            .lcout(M_this_ext_address_qZ0Z_9),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_8),
            .carryout(un1_M_this_ext_address_q_cry_9),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_10_LC_21_25_2.C_ON=1'b1;
    defparam M_this_ext_address_q_10_LC_21_25_2.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_10_LC_21_25_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_10_LC_21_25_2 (
            .in0(N__37632),
            .in1(N__37083),
            .in2(N__37243),
            .in3(N__37226),
            .lcout(M_this_ext_address_qZ0Z_10),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_9),
            .carryout(un1_M_this_ext_address_q_cry_10),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_11_LC_21_25_3.C_ON=1'b1;
    defparam M_this_ext_address_q_11_LC_21_25_3.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_11_LC_21_25_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_11_LC_21_25_3 (
            .in0(N__37874),
            .in1(N__37087),
            .in2(N__37210),
            .in3(N__37193),
            .lcout(M_this_ext_address_qZ0Z_11),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_10),
            .carryout(un1_M_this_ext_address_q_cry_11),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_12_LC_21_25_4.C_ON=1'b1;
    defparam M_this_ext_address_q_12_LC_21_25_4.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_12_LC_21_25_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_12_LC_21_25_4 (
            .in0(N__37499),
            .in1(N__37084),
            .in2(N__37180),
            .in3(N__37163),
            .lcout(M_this_ext_address_qZ0Z_12),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_11),
            .carryout(un1_M_this_ext_address_q_cry_12),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_13_LC_21_25_5.C_ON=1'b1;
    defparam M_this_ext_address_q_13_LC_21_25_5.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_13_LC_21_25_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_13_LC_21_25_5 (
            .in0(N__38903),
            .in1(N__37088),
            .in2(N__37150),
            .in3(N__37133),
            .lcout(M_this_ext_address_qZ0Z_13),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_12),
            .carryout(un1_M_this_ext_address_q_cry_13),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_14_LC_21_25_6.C_ON=1'b1;
    defparam M_this_ext_address_q_14_LC_21_25_6.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_14_LC_21_25_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 M_this_ext_address_q_14_LC_21_25_6 (
            .in0(N__37340),
            .in1(N__37085),
            .in2(N__37117),
            .in3(N__37100),
            .lcout(M_this_ext_address_qZ0Z_14),
            .ltout(),
            .carryin(un1_M_this_ext_address_q_cry_13),
            .carryout(un1_M_this_ext_address_q_cry_14),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam M_this_ext_address_q_15_LC_21_25_7.C_ON=1'b0;
    defparam M_this_ext_address_q_15_LC_21_25_7.SEQ_MODE=4'b1000;
    defparam M_this_ext_address_q_15_LC_21_25_7.LUT_INIT=16'b1101000111100010;
    LogicCell40 M_this_ext_address_q_15_LC_21_25_7 (
            .in0(N__37003),
            .in1(N__37089),
            .in2(N__38773),
            .in3(N__37022),
            .lcout(M_this_ext_address_qZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39403),
            .ce(),
            .sr(N__36818));
    defparam \this_start_data_delay.M_last_q_RNIO2A13_LC_22_20_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIO2A13_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIO2A13_LC_22_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \this_start_data_delay.M_last_q_RNIO2A13_LC_22_20_1  (
            .in0(N__36629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38346),
            .lcout(\this_start_data_delay.N_231_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIJ68N1_LC_22_20_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIJ68N1_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIJ68N1_LC_22_20_4 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \this_start_data_delay.M_last_q_RNIJ68N1_LC_22_20_4  (
            .in0(N__36951),
            .in1(N__36591),
            .in2(N__36422),
            .in3(N__36630),
            .lcout(),
            .ltout(\this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_state_q_10_LC_22_20_5.C_ON=1'b0;
    defparam M_this_state_q_10_LC_22_20_5.SEQ_MODE=4'b1000;
    defparam M_this_state_q_10_LC_22_20_5.LUT_INIT=16'b0111000000100000;
    LogicCell40 M_this_state_q_10_LC_22_20_5 (
            .in0(N__36592),
            .in1(N__38347),
            .in2(N__36575),
            .in3(N__36543),
            .lcout(M_this_state_qZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39378),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_a2_1_7_LC_22_22_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_a2_1_7_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_this_state_q_srsts_i_i_a2_1_7_LC_22_22_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \this_start_data_delay.M_this_state_q_srsts_i_i_a2_1_7_LC_22_22_0  (
            .in0(N__38343),
            .in1(N__38283),
            .in2(_gnd_net_),
            .in3(N__38164),
            .lcout(\this_start_data_delay.N_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_22_25_0 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_22_25_0 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI497F1_LC_22_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI497F1_LC_22_25_0  (
            .in0(N__38127),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38620),
            .lcout(M_this_map_ram_write_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam led_1_7_6__m7_0_a4_0_a2_0_a2_LC_23_18_0.C_ON=1'b0;
    defparam led_1_7_6__m7_0_a4_0_a2_0_a2_LC_23_18_0.SEQ_MODE=4'b0000;
    defparam led_1_7_6__m7_0_a4_0_a2_0_a2_LC_23_18_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 led_1_7_6__m7_0_a4_0_a2_0_a2_LC_23_18_0 (
            .in0(_gnd_net_),
            .in1(N__38008),
            .in2(_gnd_net_),
            .in3(N__37943),
            .lcout(led_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_24_24_1 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_24_24_1 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI7C7F1_LC_24_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI7C7F1_LC_24_24_1  (
            .in0(N__37861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38624),
            .lcout(M_this_map_ram_write_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_24_25_2 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_24_25_2 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI5A7F1_LC_24_25_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI5A7F1_LC_24_25_2  (
            .in0(N__37752),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38626),
            .lcout(M_this_map_ram_write_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_24_25_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_24_25_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI6B7F1_LC_24_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI6B7F1_LC_24_25_3  (
            .in0(N__38627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37611),
            .lcout(M_this_map_ram_write_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_24_25_5 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_24_25_5 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI8D7F1_LC_24_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI8D7F1_LC_24_25_5  (
            .in0(N__38628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37475),
            .lcout(M_this_map_ram_write_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_24_25_7 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_24_25_7 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIAF7F1_LC_24_25_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIAF7F1_LC_24_25_7  (
            .in0(N__38629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37312),
            .lcout(M_this_map_ram_write_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_24_27_3 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_24_27_3 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNI9E7F1_LC_24_27_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNI9E7F1_LC_24_27_3  (
            .in0(N__38886),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38618),
            .lcout(M_this_map_ram_write_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_24_27_4 .C_ON=1'b0;
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_24_27_4 .SEQ_MODE=4'b0000;
    defparam \this_start_data_delay.M_last_q_RNIBG7F1_LC_24_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \this_start_data_delay.M_last_q_RNIBG7F1_LC_24_27_4  (
            .in0(N__38619),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38774),
            .lcout(M_this_map_ram_write_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam M_this_map_address_q_0_LC_26_25_0.C_ON=1'b1;
    defparam M_this_map_address_q_0_LC_26_25_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_0_LC_26_25_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_0_LC_26_25_0 (
            .in0(N__39517),
            .in1(N__38509),
            .in2(N__38602),
            .in3(N__38587),
            .lcout(M_this_map_address_qZ0Z_0),
            .ltout(),
            .carryin(bfn_26_25_0_),
            .carryout(un1_M_this_map_address_q_cry_0),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_1_LC_26_25_1.C_ON=1'b1;
    defparam M_this_map_address_q_1_LC_26_25_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_1_LC_26_25_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_1_LC_26_25_1 (
            .in0(N__39523),
            .in1(N__38479),
            .in2(_gnd_net_),
            .in3(N__38465),
            .lcout(M_this_map_address_qZ0Z_1),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_0),
            .carryout(un1_M_this_map_address_q_cry_1),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_2_LC_26_25_2.C_ON=1'b1;
    defparam M_this_map_address_q_2_LC_26_25_2.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_2_LC_26_25_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_2_LC_26_25_2 (
            .in0(N__39518),
            .in1(N__38449),
            .in2(_gnd_net_),
            .in3(N__38435),
            .lcout(M_this_map_address_qZ0Z_2),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_1),
            .carryout(un1_M_this_map_address_q_cry_2),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_3_LC_26_25_3.C_ON=1'b1;
    defparam M_this_map_address_q_3_LC_26_25_3.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_3_LC_26_25_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_3_LC_26_25_3 (
            .in0(N__39524),
            .in1(N__38422),
            .in2(_gnd_net_),
            .in3(N__38408),
            .lcout(M_this_map_address_qZ0Z_3),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_2),
            .carryout(un1_M_this_map_address_q_cry_3),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_4_LC_26_25_4.C_ON=1'b1;
    defparam M_this_map_address_q_4_LC_26_25_4.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_4_LC_26_25_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_4_LC_26_25_4 (
            .in0(N__39519),
            .in1(N__38392),
            .in2(_gnd_net_),
            .in3(N__38378),
            .lcout(M_this_map_address_qZ0Z_4),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_3),
            .carryout(un1_M_this_map_address_q_cry_4),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_5_LC_26_25_5.C_ON=1'b1;
    defparam M_this_map_address_q_5_LC_26_25_5.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_5_LC_26_25_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_5_LC_26_25_5 (
            .in0(N__39521),
            .in1(N__38365),
            .in2(_gnd_net_),
            .in3(N__38351),
            .lcout(M_this_map_address_qZ0Z_5),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_4),
            .carryout(un1_M_this_map_address_q_cry_5),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_6_LC_26_25_6.C_ON=1'b1;
    defparam M_this_map_address_q_6_LC_26_25_6.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_6_LC_26_25_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_6_LC_26_25_6 (
            .in0(N__39520),
            .in1(N__39607),
            .in2(_gnd_net_),
            .in3(N__39593),
            .lcout(M_this_map_address_qZ0Z_6),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_5),
            .carryout(un1_M_this_map_address_q_cry_6),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_7_LC_26_25_7.C_ON=1'b1;
    defparam M_this_map_address_q_7_LC_26_25_7.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_7_LC_26_25_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_7_LC_26_25_7 (
            .in0(N__39522),
            .in1(N__39577),
            .in2(_gnd_net_),
            .in3(N__39563),
            .lcout(M_this_map_address_qZ0Z_7),
            .ltout(),
            .carryin(un1_M_this_map_address_q_cry_6),
            .carryout(un1_M_this_map_address_q_cry_7),
            .clk(N__39424),
            .ce(),
            .sr(N__38956));
    defparam M_this_map_address_q_8_LC_26_26_0.C_ON=1'b1;
    defparam M_this_map_address_q_8_LC_26_26_0.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_8_LC_26_26_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 M_this_map_address_q_8_LC_26_26_0 (
            .in0(N__39525),
            .in1(N__39547),
            .in2(_gnd_net_),
            .in3(N__39533),
            .lcout(M_this_map_address_qZ0Z_8),
            .ltout(),
            .carryin(bfn_26_26_0_),
            .carryout(un1_M_this_map_address_q_cry_8),
            .clk(N__39430),
            .ce(),
            .sr(N__38955));
    defparam M_this_map_address_q_9_LC_26_26_1.C_ON=1'b0;
    defparam M_this_map_address_q_9_LC_26_26_1.SEQ_MODE=4'b1000;
    defparam M_this_map_address_q_9_LC_26_26_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 M_this_map_address_q_9_LC_26_26_1 (
            .in0(N__39448),
            .in1(N__39526),
            .in2(_gnd_net_),
            .in3(N__39464),
            .lcout(M_this_map_address_qZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__39430),
            .ce(),
            .sr(N__38955));
endmodule // cu_top_0
