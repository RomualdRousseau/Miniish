-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec 10 2020 17:47:04

-- File Generated:     Jun 1 2022 00:08:23

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cu_top_0" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cu_top_0
entity cu_top_0 is
port (
    port_address : inout std_logic_vector(15 downto 0);
    port_data : in std_logic_vector(7 downto 0);
    debug : out std_logic_vector(1 downto 0);
    rgb : out std_logic_vector(5 downto 0);
    led : out std_logic_vector(7 downto 0);
    vsync : out std_logic;
    vblank : out std_logic;
    rst_n : in std_logic;
    port_rw : inout std_logic;
    port_nmib : out std_logic;
    port_enb : in std_logic;
    port_dmab : out std_logic;
    port_data_rw : out std_logic;
    port_clk : in std_logic;
    hsync : out std_logic;
    hblank : out std_logic;
    clk : in std_logic);
end cu_top_0;

-- Architecture of cu_top_0
-- View name is \INTERFACE\
architecture \INTERFACE\ of cu_top_0 is

signal \N__40097\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40086\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40084\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40076\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40068\ : std_logic;
signal \N__40067\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40058\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40049\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40040\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40032\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40023\ : std_logic;
signal \N__40022\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40013\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40004\ : std_logic;
signal \N__40003\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39995\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39968\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39959\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39950\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39941\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39932\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39923\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39914\ : std_logic;
signal \N__39913\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39904\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39896\ : std_logic;
signal \N__39895\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39886\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39877\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39868\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39851\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39806\ : std_logic;
signal \N__39805\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39788\ : std_logic;
signal \N__39787\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39778\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39769\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39760\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39752\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39734\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39716\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39698\ : std_logic;
signal \N__39697\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39688\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39661\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39652\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39644\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39635\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39593\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39577\ : std_logic;
signal \N__39574\ : std_logic;
signal \N__39571\ : std_logic;
signal \N__39568\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39544\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39530\ : std_logic;
signal \N__39527\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39524\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39519\ : std_logic;
signal \N__39518\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39491\ : std_logic;
signal \N__39488\ : std_logic;
signal \N__39481\ : std_logic;
signal \N__39478\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39472\ : std_logic;
signal \N__39469\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39432\ : std_logic;
signal \N__39431\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39428\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39419\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39416\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39413\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39410\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39407\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39404\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39398\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39395\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39388\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39385\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39380\ : std_logic;
signal \N__39379\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39377\ : std_logic;
signal \N__39376\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39368\ : std_logic;
signal \N__39367\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39364\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39361\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39358\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39355\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39348\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39342\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39339\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39335\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39333\ : std_logic;
signal \N__39332\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39320\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39312\ : std_logic;
signal \N__39311\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39302\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39299\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39294\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39291\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39284\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__38969\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38963\ : std_logic;
signal \N__38962\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38956\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38953\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38951\ : std_logic;
signal \N__38924\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38918\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38911\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38890\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38839\ : std_logic;
signal \N__38836\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38801\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38780\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38765\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38738\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38655\ : std_logic;
signal \N__38652\ : std_logic;
signal \N__38649\ : std_logic;
signal \N__38646\ : std_logic;
signal \N__38641\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38633\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38629\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38559\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38513\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38483\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38465\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38440\ : std_logic;
signal \N__38435\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38399\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38392\ : std_logic;
signal \N__38389\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38378\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38362\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38351\ : std_logic;
signal \N__38348\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38284\ : std_logic;
signal \N__38283\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38281\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38274\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38258\ : std_logic;
signal \N__38255\ : std_logic;
signal \N__38252\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38180\ : std_logic;
signal \N__38171\ : std_logic;
signal \N__38168\ : std_logic;
signal \N__38165\ : std_logic;
signal \N__38164\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38141\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38135\ : std_logic;
signal \N__38132\ : std_logic;
signal \N__38129\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38102\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38093\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38069\ : std_logic;
signal \N__38066\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38042\ : std_logic;
signal \N__38039\ : std_logic;
signal \N__38036\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38024\ : std_logic;
signal \N__38021\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38015\ : std_logic;
signal \N__38012\ : std_logic;
signal \N__38009\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37997\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37993\ : std_logic;
signal \N__37990\ : std_logic;
signal \N__37987\ : std_logic;
signal \N__37984\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37979\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37961\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37943\ : std_logic;
signal \N__37940\ : std_logic;
signal \N__37939\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37907\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37892\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37861\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37853\ : std_logic;
signal \N__37852\ : std_logic;
signal \N__37847\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37756\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37751\ : std_logic;
signal \N__37746\ : std_logic;
signal \N__37743\ : std_logic;
signal \N__37740\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37735\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37668\ : std_logic;
signal \N__37665\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37637\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37615\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37579\ : std_logic;
signal \N__37576\ : std_logic;
signal \N__37571\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37560\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37535\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37523\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37517\ : std_logic;
signal \N__37514\ : std_logic;
signal \N__37511\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37499\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37493\ : std_logic;
signal \N__37490\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37472\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37466\ : std_logic;
signal \N__37463\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37435\ : std_logic;
signal \N__37432\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37406\ : std_logic;
signal \N__37403\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37393\ : std_logic;
signal \N__37390\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37382\ : std_logic;
signal \N__37379\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37375\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37352\ : std_logic;
signal \N__37351\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37331\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37312\ : std_logic;
signal \N__37309\ : std_logic;
signal \N__37306\ : std_logic;
signal \N__37303\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37292\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37286\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37280\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37267\ : std_logic;
signal \N__37264\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37256\ : std_logic;
signal \N__37253\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37243\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37234\ : std_logic;
signal \N__37231\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37223\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37210\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37201\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37193\ : std_logic;
signal \N__37190\ : std_logic;
signal \N__37187\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37181\ : std_logic;
signal \N__37180\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37157\ : std_logic;
signal \N__37154\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37133\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37124\ : std_logic;
signal \N__37121\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37105\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37094\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37085\ : std_logic;
signal \N__37084\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37033\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37022\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36970\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36962\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36943\ : std_logic;
signal \N__36940\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36906\ : std_logic;
signal \N__36903\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36887\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36845\ : std_logic;
signal \N__36844\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36841\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36835\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36832\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36829\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36809\ : std_logic;
signal \N__36806\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36776\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36580\ : std_logic;
signal \N__36575\ : std_logic;
signal \N__36572\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36566\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36521\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36515\ : std_logic;
signal \N__36512\ : std_logic;
signal \N__36509\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36448\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36421\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36392\ : std_logic;
signal \N__36389\ : std_logic;
signal \N__36386\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36344\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36338\ : std_logic;
signal \N__36335\ : std_logic;
signal \N__36332\ : std_logic;
signal \N__36329\ : std_logic;
signal \N__36328\ : std_logic;
signal \N__36325\ : std_logic;
signal \N__36322\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36308\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36301\ : std_logic;
signal \N__36298\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36281\ : std_logic;
signal \N__36278\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36257\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36251\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36200\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36178\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36170\ : std_logic;
signal \N__36167\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36160\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36122\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36097\ : std_logic;
signal \N__36094\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36034\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36008\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35980\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35962\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35945\ : std_logic;
signal \N__35942\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35914\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35851\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35809\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35712\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35612\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35599\ : std_logic;
signal \N__35596\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35585\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35536\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35460\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35437\ : std_logic;
signal \N__35434\ : std_logic;
signal \N__35431\ : std_logic;
signal \N__35426\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35336\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35246\ : std_logic;
signal \N__35243\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35186\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35141\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35072\ : std_logic;
signal \N__35069\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35055\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35006\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34993\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34954\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34862\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34829\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34824\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34757\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34703\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34672\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34658\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34649\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34519\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34510\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34484\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34448\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34432\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34394\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34388\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34379\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34352\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34235\ : std_logic;
signal \N__34232\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34226\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34178\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34088\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34079\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34069\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34019\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34016\ : std_logic;
signal \N__34013\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33913\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33767\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33742\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33664\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33646\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33632\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33620\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33611\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33599\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33572\ : std_logic;
signal \N__33569\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33536\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33532\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33477\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33467\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33410\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33407\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33385\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33272\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33250\ : std_logic;
signal \N__33245\ : std_logic;
signal \N__33242\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33212\ : std_logic;
signal \N__33209\ : std_logic;
signal \N__33206\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33200\ : std_logic;
signal \N__33197\ : std_logic;
signal \N__33194\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33131\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33092\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33074\ : std_logic;
signal \N__33071\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33029\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32708\ : std_logic;
signal \N__32705\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32627\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32584\ : std_logic;
signal \N__32581\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32564\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32562\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32544\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32514\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32492\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32411\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32324\ : std_logic;
signal \N__32321\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32264\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32210\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32195\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32189\ : std_logic;
signal \N__32186\ : std_logic;
signal \N__32183\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32126\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32107\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31898\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31889\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31838\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31819\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31738\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31735\ : std_logic;
signal \N__31732\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31711\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31693\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31675\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31661\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31598\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31496\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31423\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31399\ : std_logic;
signal \N__31396\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31316\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31286\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31274\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31187\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31175\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31136\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31130\ : std_logic;
signal \N__31129\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31034\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30954\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30802\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30757\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30719\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30689\ : std_logic;
signal \N__30686\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30674\ : std_logic;
signal \N__30671\ : std_logic;
signal \N__30668\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30656\ : std_logic;
signal \N__30653\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30635\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30599\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30572\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30545\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30509\ : std_logic;
signal \N__30506\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30326\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30282\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30254\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30236\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30221\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30167\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30152\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29903\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29795\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29770\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29602\ : std_logic;
signal \N__29599\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29551\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29494\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29302\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29290\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29255\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29085\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28972\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28891\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28742\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28466\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28444\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28346\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28223\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28006\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27968\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27932\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27882\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27839\ : std_logic;
signal \N__27836\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27497\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27434\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27320\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27197\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26684\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25798\ : std_logic;
signal \N__25797\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25661\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25070\ : std_logic;
signal \N__25067\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24853\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24614\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24253\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24209\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23558\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23317\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19598\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15071\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal port_data_rw_0_i : std_logic;
signal port_clk_c : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_0\ : std_logic;
signal rgb_c_3 : std_logic;
signal rgb_c_1 : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_1\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_2\ : std_logic;
signal rgb_c_2 : std_logic;
signal rgb_c_4 : std_logic;
signal rgb_c_5 : std_logic;
signal \M_this_vga_signals_address_6\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_cascade_\ : std_logic;
signal \M_this_vga_signals_address_1\ : std_logic;
signal \this_vga_signals.SUM_3_1\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_axbxc3_1_2\ : std_logic;
signal \this_vga_signals.un2_hsynclto6_0\ : std_logic;
signal \this_vga_signals.un4_hsynclt7_cascade_\ : std_logic;
signal \this_vga_signals.hsync_1_1\ : std_logic;
signal \this_vga_signals.un4_hsynclt8_0_cascade_\ : std_logic;
signal this_vga_signals_hsync_1_i : std_logic;
signal this_vga_signals_hvisibility_i : std_logic;
signal this_vga_signals_vvisibility_i : std_logic;
signal rgb_c_0 : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3\ : std_logic;
signal \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \M_this_vga_signals_address_2\ : std_logic;
signal \this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_\ : std_logic;
signal \this_vga_signals.if_m7_0_o4_1_ns_1\ : std_logic;
signal \this_vga_signals.SUM_3_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.mult1_un89_sum_c3_0\ : std_logic;
signal \M_this_vga_signals_address_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_2\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_2_cascade_\ : std_logic;
signal \M_this_vga_signals_address_3\ : std_logic;
signal \M_this_vga_signals_address_5\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axbxc3_2\ : std_logic;
signal \M_this_vga_signals_address_4\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\ : std_logic;
signal \this_vga_signals.SUM_3\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m1_1\ : std_logic;
signal \this_vga_ramdac.N_3139_reto\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_7\ : std_logic;
signal \this_vga_signals.un1_M_hcounter_d_cry_8\ : std_logic;
signal \bfn_7_18_0_\ : std_logic;
signal \M_this_oam_ram_read_data_14\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_14\ : std_logic;
signal \M_this_oam_ram_read_data_15\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_15\ : std_logic;
signal \this_ppu.oam_cache.N_823_0\ : std_logic;
signal \this_ppu.oam_cache.N_820_0\ : std_logic;
signal \M_this_oam_ram_read_data_8\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_8\ : std_logic;
signal \M_this_oam_ram_read_data_9\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_9\ : std_logic;
signal \M_this_oam_ram_read_data_10\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_10\ : std_logic;
signal \bfn_7_20_0_\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_3\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_4\ : std_logic;
signal \this_ppu.m71_i_o2_0_cascade_\ : std_logic;
signal \this_ppu.m71_i_o2_1\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_0\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_qZ0Z_3\ : std_logic;
signal \this_ppu.oam_cache.N_826_0\ : std_logic;
signal \this_ppu.oam_cache.N_824_0\ : std_logic;
signal \this_ppu.oam_cache.N_821_0\ : std_logic;
signal \this_ppu.oam_cache.N_822_0\ : std_logic;
signal \this_ppu.oam_cache.N_819_0\ : std_logic;
signal \this_ppu.oam_cache.N_825_0\ : std_logic;
signal \M_this_oam_ram_read_data_0\ : std_logic;
signal \M_this_oam_ram_read_data_6\ : std_logic;
signal \M_this_oam_ram_read_data_1\ : std_logic;
signal \M_this_oam_ram_read_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_7\ : std_logic;
signal \M_this_oam_ram_read_data_4\ : std_logic;
signal \M_this_oam_ram_read_data_5\ : std_logic;
signal \M_this_oam_ram_read_data_2\ : std_logic;
signal \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_\ : std_logic;
signal \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4\ : std_logic;
signal \this_ppu.m35_i_a2_3_cascade_\ : std_logic;
signal \this_ppu.N_802_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_1\ : std_logic;
signal \this_vga_signals.un2_hsynclto3_1_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_4\ : std_logic;
signal \this_vga_ramdac.M_this_vga_ramdac_en_reto\ : std_logic;
signal \this_vga_ramdac.i2_mux_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3140_reto\ : std_logic;
signal \this_vga_ramdac.N_24_mux_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3138_reto\ : std_logic;
signal \this_ppu.oam_cache.mem_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.M_hcounter_d7lt7_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_6\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_8\ : std_logic;
signal \this_vga_signals.N_864_cascade_\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_7\ : std_logic;
signal \this_vga_ramdac.m16_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3141_reto\ : std_logic;
signal \this_vga_ramdac.m19_cascade_\ : std_logic;
signal \this_vga_ramdac.N_3142_reto\ : std_logic;
signal \M_this_vram_read_data_0\ : std_logic;
signal \M_this_vram_read_data_2\ : std_logic;
signal \M_this_vram_read_data_3\ : std_logic;
signal \M_this_vram_read_data_1\ : std_logic;
signal \this_vga_ramdac.m6\ : std_logic;
signal \this_ppu.oam_cache.mem_17\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_17\ : std_logic;
signal \this_ppu.oam_cache.mem_16\ : std_logic;
signal \this_vga_ramdac.i2_mux_0\ : std_logic;
signal \this_vga_ramdac.N_3143_reto\ : std_logic;
signal \this_ppu.oam_cache.mem_18\ : std_logic;
signal \this_ppu.N_777_0\ : std_logic;
signal \this_ppu.N_776_0\ : std_logic;
signal \this_ppu.N_932_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_state_q_7_i_0_0_cascade_\ : std_logic;
signal \this_ppu.N_775_0\ : std_logic;
signal \this_ppu.N_932_0\ : std_logic;
signal \this_ppu.N_838_7\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_16\ : std_logic;
signal \bfn_9_21_0_\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_17\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_0\ : std_logic;
signal \this_ppu.M_this_oam_ram_read_data_i_18\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_1\ : std_logic;
signal \this_ppu.m28_e_i_o2_0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_2\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_3\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_4\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_5\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_6\ : std_logic;
signal \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_21\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_22\ : std_logic;
signal \M_this_oam_ram_read_data_i_22\ : std_logic;
signal \M_this_oam_ram_read_data_23\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_23\ : std_logic;
signal \M_this_oam_ram_read_data_24\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_24\ : std_logic;
signal \M_this_oam_ram_read_data_25\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_25\ : std_logic;
signal \M_this_oam_ram_read_data_26\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_26\ : std_logic;
signal \M_this_oam_ram_write_data_14\ : std_logic;
signal \M_this_oam_ram_read_data_30\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_30\ : std_logic;
signal \M_this_oam_ram_write_data_13\ : std_logic;
signal \M_this_oam_ram_write_data_15\ : std_logic;
signal \M_this_oam_ram_write_data_18\ : std_logic;
signal \M_this_oam_ram_read_data_31\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_31\ : std_logic;
signal \M_this_oam_ram_write_data_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_3\ : std_logic;
signal \M_this_oam_ram_write_data_3\ : std_logic;
signal \M_this_oam_ram_read_data_21\ : std_logic;
signal \M_this_oam_ram_read_data_i_21\ : std_logic;
signal \M_this_data_tmp_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_write_data_6\ : std_logic;
signal \M_this_oam_ram_write_data_5\ : std_logic;
signal \M_this_oam_ram_write_data_7\ : std_logic;
signal \M_this_oam_ram_read_data_28\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_28\ : std_logic;
signal \M_this_oam_ram_read_data_29\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_29\ : std_logic;
signal \M_this_oam_ram_write_data_16\ : std_logic;
signal \M_this_oam_ram_write_data_22\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_19\ : std_logic;
signal \M_this_oam_ram_read_data_i_19\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_20\ : std_logic;
signal \M_this_oam_ram_read_data_i_20\ : std_logic;
signal \M_this_oam_ram_write_data_27\ : std_logic;
signal \M_this_oam_ram_write_data_30\ : std_logic;
signal \M_this_oam_ram_write_data_17\ : std_logic;
signal \M_this_oam_ram_write_data_29\ : std_logic;
signal \M_this_oam_ram_write_data_24\ : std_logic;
signal dma_0_i : std_logic;
signal \this_ppu.oam_cache.mem_7\ : std_logic;
signal \this_ppu.oam_cache.mem_3\ : std_logic;
signal \this_ppu.oam_cache.mem_4\ : std_logic;
signal \this_pixel_clk_M_counter_q_i_1\ : std_logic;
signal \this_pixel_clk_M_counter_q_0\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_hcounter_qZ0Z_0\ : std_logic;
signal \N_3_0_cascade_\ : std_logic;
signal \this_vga_signals.M_pcounter_q_i_2_0\ : std_logic;
signal \this_vga_signals.M_pcounter_q_3_0\ : std_logic;
signal \this_vga_signals.N_1188_1\ : std_logic;
signal \this_vga_signals.N_1188_1_cascade_\ : std_logic;
signal \this_vga_signals.N_933_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_pcounter_qZ0Z_0\ : std_logic;
signal \N_2_0\ : std_logic;
signal \M_this_vga_signals_pixel_clk_0_0\ : std_logic;
signal \N_2_0_cascade_\ : std_logic;
signal \N_3_0\ : std_logic;
signal \G_462\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_16\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_17\ : std_logic;
signal \M_this_ppu_spr_addr_4\ : std_logic;
signal \this_ppu.offset_y_cry_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_18\ : std_logic;
signal \this_ppu.offset_y_cry_1\ : std_logic;
signal \M_this_ppu_spr_addr_5\ : std_logic;
signal \this_ppu.oam_cache.mem_10\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_10\ : std_logic;
signal \this_ppu.N_836_cascade_\ : std_logic;
signal \this_ppu.oam_cache.mem_9\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_2\ : std_logic;
signal \un1_M_this_warmup_d_cry_1\ : std_logic;
signal \M_this_warmup_qZ0Z_3\ : std_logic;
signal \un1_M_this_warmup_d_cry_2\ : std_logic;
signal \M_this_warmup_qZ0Z_4\ : std_logic;
signal \un1_M_this_warmup_d_cry_3\ : std_logic;
signal \M_this_warmup_qZ0Z_5\ : std_logic;
signal \un1_M_this_warmup_d_cry_4\ : std_logic;
signal \M_this_warmup_qZ0Z_6\ : std_logic;
signal \un1_M_this_warmup_d_cry_5\ : std_logic;
signal \M_this_warmup_qZ0Z_7\ : std_logic;
signal \un1_M_this_warmup_d_cry_6\ : std_logic;
signal \M_this_warmup_qZ0Z_8\ : std_logic;
signal \un1_M_this_warmup_d_cry_7\ : std_logic;
signal \un1_M_this_warmup_d_cry_8\ : std_logic;
signal \M_this_warmup_qZ0Z_9\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_10\ : std_logic;
signal \un1_M_this_warmup_d_cry_9\ : std_logic;
signal \M_this_warmup_qZ0Z_11\ : std_logic;
signal \un1_M_this_warmup_d_cry_10\ : std_logic;
signal \M_this_warmup_qZ0Z_12\ : std_logic;
signal \un1_M_this_warmup_d_cry_11\ : std_logic;
signal \M_this_warmup_qZ0Z_13\ : std_logic;
signal \un1_M_this_warmup_d_cry_12\ : std_logic;
signal \M_this_warmup_qZ0Z_14\ : std_logic;
signal \un1_M_this_warmup_d_cry_13\ : std_logic;
signal \M_this_warmup_qZ0Z_15\ : std_logic;
signal \un1_M_this_warmup_d_cry_14\ : std_logic;
signal \M_this_warmup_qZ0Z_16\ : std_logic;
signal \un1_M_this_warmup_d_cry_15\ : std_logic;
signal \un1_M_this_warmup_d_cry_16\ : std_logic;
signal \M_this_warmup_qZ0Z_17\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_18\ : std_logic;
signal \un1_M_this_warmup_d_cry_17\ : std_logic;
signal \M_this_warmup_qZ0Z_19\ : std_logic;
signal \un1_M_this_warmup_d_cry_18\ : std_logic;
signal \M_this_warmup_qZ0Z_20\ : std_logic;
signal \un1_M_this_warmup_d_cry_19\ : std_logic;
signal \M_this_warmup_qZ0Z_21\ : std_logic;
signal \un1_M_this_warmup_d_cry_20\ : std_logic;
signal \M_this_warmup_qZ0Z_22\ : std_logic;
signal \un1_M_this_warmup_d_cry_21\ : std_logic;
signal \M_this_warmup_qZ0Z_23\ : std_logic;
signal \un1_M_this_warmup_d_cry_22\ : std_logic;
signal \M_this_warmup_qZ0Z_24\ : std_logic;
signal \un1_M_this_warmup_d_cry_23\ : std_logic;
signal \un1_M_this_warmup_d_cry_24\ : std_logic;
signal \M_this_warmup_qZ0Z_25\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \M_this_warmup_qZ0Z_26\ : std_logic;
signal \un1_M_this_warmup_d_cry_25\ : std_logic;
signal \M_this_warmup_qZ0Z_27\ : std_logic;
signal \un1_M_this_warmup_d_cry_26\ : std_logic;
signal \un1_M_this_warmup_d_cry_27\ : std_logic;
signal \M_this_warmup_qZ0Z_28\ : std_logic;
signal \M_this_data_tmp_qZ0Z_8\ : std_logic;
signal \M_this_data_tmp_qZ0Z_14\ : std_logic;
signal \M_this_data_tmp_qZ0Z_10\ : std_logic;
signal \M_this_oam_ram_write_data_10\ : std_logic;
signal \M_this_oam_ram_write_data_12\ : std_logic;
signal \M_this_data_tmp_qZ0Z_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_5\ : std_logic;
signal \M_this_data_tmp_qZ0Z_22\ : std_logic;
signal \M_this_data_tmp_qZ0Z_16\ : std_logic;
signal \M_this_oam_ram_write_data_31\ : std_logic;
signal \M_this_oam_ram_write_data_21\ : std_logic;
signal \M_this_oam_ram_write_data_23\ : std_logic;
signal \this_spr_ram.mem_WE_12\ : std_logic;
signal \this_spr_ram.mem_WE_14\ : std_logic;
signal \this_ppu.oam_cache.mem_5\ : std_logic;
signal \this_spr_ram.mem_WE_0\ : std_logic;
signal \N_34_i\ : std_logic;
signal \this_ppu.oam_cache.mem_14\ : std_logic;
signal \this_ppu.M_oam_curr_qc_0_1_cascade_\ : std_logic;
signal \this_ppu.m35_i_a2_4\ : std_logic;
signal \this_ppu.N_827_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c5\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c5_cascade_\ : std_logic;
signal \M_this_ppu_vram_addr_5\ : std_logic;
signal \M_this_ppu_vram_addr_6\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c2\ : std_logic;
signal \M_this_ppu_vram_addr_1\ : std_logic;
signal \M_this_ppu_vram_addr_0\ : std_logic;
signal \M_this_ppu_vram_addr_2\ : std_logic;
signal \this_ppu.N_827_0\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c3_cascade_\ : std_logic;
signal \M_this_ppu_vram_addr_4\ : std_logic;
signal \this_ppu.N_1210_0\ : std_logic;
signal \this_ppu.un1_M_screen_x_q_c3\ : std_logic;
signal \this_ppu.oam_cache.mem_13\ : std_logic;
signal \this_ppu.oam_cache.mem_12\ : std_logic;
signal \this_ppu.m13_0_a2_0_0\ : std_logic;
signal \this_ppu.N_844_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_1\ : std_logic;
signal \M_this_warmup_qZ0Z_1\ : std_logic;
signal \M_this_warmup_qZ0Z_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_9\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_16\ : std_logic;
signal \M_this_ppu_spr_addr_3\ : std_logic;
signal \this_ppu.M_state_qZ0Z_2\ : std_logic;
signal \M_this_oam_address_qZ0Z_6\ : std_logic;
signal \M_this_oam_address_qZ0Z_7\ : std_logic;
signal \M_this_data_tmp_qZ0Z_12\ : std_logic;
signal \M_this_data_tmp_qZ0Z_15\ : std_logic;
signal \M_this_data_tmp_qZ0Z_13\ : std_logic;
signal \M_this_oam_ram_write_data_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_20\ : std_logic;
signal \M_this_oam_ram_write_data_20\ : std_logic;
signal \M_this_oam_ram_write_data_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_9\ : std_logic;
signal \M_this_oam_ram_write_data_9\ : std_logic;
signal \M_this_oam_ram_write_data_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_11\ : std_logic;
signal \M_this_oam_ram_write_data_11\ : std_logic;
signal \M_this_data_tmp_qZ0Z_17\ : std_logic;
signal \M_this_data_tmp_qZ0Z_23\ : std_logic;
signal \M_this_oam_ram_write_data_19\ : std_logic;
signal \M_this_oam_ram_write_data_28\ : std_logic;
signal \M_this_oam_ram_write_data_25\ : std_logic;
signal \this_spr_ram.mem_out_bus4_1\ : std_logic;
signal \this_spr_ram.mem_out_bus0_1\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\ : std_logic;
signal \this_spr_ram.mem_out_bus5_1\ : std_logic;
signal \this_spr_ram.mem_out_bus1_1\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus7_1\ : std_logic;
signal \this_spr_ram.mem_out_bus3_1\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus6_1\ : std_logic;
signal \this_spr_ram.mem_out_bus2_1\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\ : std_logic;
signal \this_spr_ram.mem_out_bus4_3\ : std_logic;
signal \this_spr_ram.mem_out_bus0_3\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\ : std_logic;
signal \M_this_ppu_vram_addr_3\ : std_logic;
signal \this_vga_signals.N_22_0_cascade_\ : std_logic;
signal \N_856_i\ : std_logic;
signal \this_spr_ram.mem_out_bus5_3\ : std_logic;
signal \this_spr_ram.mem_out_bus1_3\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3\ : std_logic;
signal \M_this_spr_ram_read_data_3_cascade_\ : std_logic;
signal \N_25_0_i\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_14\ : std_logic;
signal \this_spr_ram.mem_out_bus4_2\ : std_logic;
signal \this_spr_ram.mem_out_bus0_2\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_6\ : std_logic;
signal \this_ppu.M_state_q_inv_1_cascade_\ : std_logic;
signal \M_this_map_ram_read_data_6\ : std_logic;
signal \this_ppu.m48_i_a2_0\ : std_logic;
signal \this_spr_ram.mem_out_bus5_2\ : std_logic;
signal \this_spr_ram.mem_out_bus1_2\ : std_logic;
signal \this_spr_ram.mem_out_bus7_2\ : std_logic;
signal \this_spr_ram.mem_out_bus3_2\ : std_logic;
signal \this_spr_ram.mem_out_bus2_2\ : std_logic;
signal \this_spr_ram.mem_out_bus6_2\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\ : std_logic;
signal \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\ : std_logic;
signal \this_ppu_N_247\ : std_logic;
signal \this_vga_signals.N_22_0\ : std_logic;
signal \M_this_spr_ram_read_data_2_cascade_\ : std_logic;
signal \N_28_0_i\ : std_logic;
signal \M_this_ppu_oam_addr_4\ : std_logic;
signal \M_this_spr_ram_read_data_2\ : std_logic;
signal \M_this_spr_ram_read_data_1\ : std_logic;
signal \M_this_spr_ram_read_data_3\ : std_logic;
signal \this_ppu.M_oam_curr_dZ0Z25_cascade_\ : std_logic;
signal \this_ppu.N_834_0\ : std_logic;
signal \M_this_ppu_oam_addr_0\ : std_logic;
signal \this_ppu.N_834_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_state_q_7_i_0_0\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c1\ : std_logic;
signal \M_this_ppu_oam_addr_1\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c1_cascade_\ : std_logic;
signal \M_this_ppu_oam_addr_2\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c3\ : std_logic;
signal \M_this_ppu_oam_addr_3\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c3_cascade_\ : std_logic;
signal \this_ppu.N_778_0\ : std_logic;
signal \this_ppu.un1_M_oam_curr_q_1_c5\ : std_logic;
signal \M_this_ppu_oam_addr_5\ : std_logic;
signal \this_ppu.M_oam_curr_qc_0_1\ : std_logic;
signal \this_ppu.M_oam_curr_qZ0Z_6\ : std_logic;
signal \M_this_status_flags_qZ0Z_0\ : std_logic;
signal \this_ppu.oam_cache.mem_15\ : std_logic;
signal \this_ppu.N_784_0\ : std_logic;
signal \this_vga_signals.N_859_cascade_\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_13\ : std_logic;
signal \this_ppu.m9_0_a2_5_cascade_\ : std_logic;
signal \this_vga_signals.i22_mux\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.M_lcounter_qZ0Z_0\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2\ : std_logic;
signal \this_ppu.N_814_cascade_\ : std_logic;
signal \this_ppu.N_806_cascade_\ : std_logic;
signal \this_ppu.N_806\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_0\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_1\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_3\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_2\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_4\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_3\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_5\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_4\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_6\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_5\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_6\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6_1Z0Z_10\ : std_logic;
signal \M_this_oam_ram_read_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_11\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6Z0Z_10\ : std_logic;
signal \M_this_oam_address_qZ0Z_3\ : std_logic;
signal \M_this_oam_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_oam_address_q_c4\ : std_logic;
signal \M_this_oam_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_oam_address_q_c4_cascade_\ : std_logic;
signal \M_this_oam_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_oam_address_q_c6\ : std_logic;
signal \N_1240_0\ : std_logic;
signal \M_this_oam_ram_write_data_0_sqmuxa_cascade_\ : std_logic;
signal \M_this_oam_ram_write_data_26\ : std_logic;
signal \M_this_oam_ram_write_data_0_sqmuxa\ : std_logic;
signal \M_this_oam_ram_write_data_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_0\ : std_logic;
signal \M_this_data_tmp_qZ0Z_4\ : std_logic;
signal \M_this_data_tmp_qZ0Z_2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_21\ : std_logic;
signal \this_spr_ram.mem_out_bus7_0\ : std_logic;
signal \this_spr_ram.mem_out_bus3_0\ : std_logic;
signal \this_spr_ram.mem_out_bus4_0\ : std_logic;
signal \this_spr_ram.mem_out_bus0_0\ : std_logic;
signal \this_spr_ram.mem_out_bus5_0\ : std_logic;
signal \this_spr_ram.mem_out_bus1_0\ : std_logic;
signal \this_spr_ram.mem_out_bus6_0\ : std_logic;
signal \this_spr_ram.mem_out_bus2_0\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_12\ : std_logic;
signal \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\ : std_logic;
signal \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\ : std_logic;
signal \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\ : std_logic;
signal \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\ : std_logic;
signal \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\ : std_logic;
signal \M_this_spr_ram_read_data_0\ : std_logic;
signal \M_this_map_ram_read_data_7\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_3\ : std_logic;
signal \M_this_map_ram_read_data_3\ : std_logic;
signal \M_this_ppu_spr_addr_9\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_4\ : std_logic;
signal \M_this_map_ram_read_data_4\ : std_logic;
signal \M_this_ppu_spr_addr_10\ : std_logic;
signal \M_this_ppu_spr_addr_0\ : std_logic;
signal \this_spr_ram.mem_out_bus6_3\ : std_logic;
signal \this_spr_ram.mem_out_bus2_3\ : std_logic;
signal \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_5\ : std_logic;
signal \M_this_map_ram_read_data_5\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_11\ : std_logic;
signal \this_ppu.N_797\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c4_cascade_\ : std_logic;
signal \this_ppu.N_802\ : std_logic;
signal \this_spr_ram.mem_out_bus7_3\ : std_logic;
signal \this_spr_ram.mem_out_bus3_3\ : std_logic;
signal \this_spr_ram.mem_radregZ0Z_13\ : std_logic;
signal \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_5\ : std_logic;
signal \this_ppu.N_796_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_8\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c6_cascade_\ : std_logic;
signal \this_ppu.N_798_0_cascade_\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c3\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c3_cascade_\ : std_logic;
signal \this_ppu.N_798_0\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c2_cascade_\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c5_cascade_\ : std_logic;
signal \this_ppu.N_800\ : std_logic;
signal \this_ppu.N_800_cascade_\ : std_logic;
signal \this_ppu.M_state_qZ0Z_11\ : std_logic;
signal \N_18\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c2\ : std_logic;
signal \this_ppu.M_oam_curr_dZ0Z25\ : std_logic;
signal \this_ppu.M_state_qZ0Z_7\ : std_logic;
signal \this_ppu.M_state_qZ0Z_9\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c1_cascade_\ : std_logic;
signal \M_this_scroll_qZ0Z_10\ : std_logic;
signal \M_this_scroll_qZ0Z_11\ : std_logic;
signal \M_this_scroll_qZ0Z_13\ : std_logic;
signal \M_this_scroll_qZ0Z_14\ : std_logic;
signal \M_this_scroll_qZ0Z_8\ : std_logic;
signal \N_829_0_cascade_\ : std_logic;
signal \N_58_0_cascade_\ : std_logic;
signal \this_ppu.N_97_mux\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_\ : std_logic;
signal \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_2\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_1\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ0Z_7\ : std_logic;
signal \this_ppu.m9_0_a2_4\ : std_logic;
signal \this_ppu.M_pixel_cnt_qZ1Z_0\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_axb_0\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6_2Z0Z_10\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6_4Z0Z_10\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6_0Z0Z_10\ : std_logic;
signal \this_ppu.M_state_qZ0Z_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_10\ : std_logic;
signal \this_ppu.N_835_0_cascade_\ : std_logic;
signal \this_ppu.N_783_cascade_\ : std_logic;
signal \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0\ : std_logic;
signal \this_ppu.oam_cache.mem_2\ : std_logic;
signal \this_ppu.N_60_0\ : std_logic;
signal \this_ppu.M_state_qZ0Z_0\ : std_logic;
signal \this_ppu.N_835_0\ : std_logic;
signal \this_ppu.N_807\ : std_logic;
signal \this_ppu.N_814\ : std_logic;
signal \this_ppu.N_783\ : std_logic;
signal \this_ppu.M_state_q_RNISP3R6_3Z0Z_10\ : std_logic;
signal \un1_M_this_oam_address_q_c2\ : std_logic;
signal \M_this_data_tmp_qZ0Z_18\ : std_logic;
signal \M_this_data_tmp_qZ0Z_1\ : std_logic;
signal \M_this_data_tmp_qZ0Z_19\ : std_logic;
signal \N_1232_0\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c6\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c4\ : std_logic;
signal \this_ppu_M_screen_y_q_3\ : std_logic;
signal \this_ppu.un3_M_screen_y_d_0_c2\ : std_logic;
signal \this_ppu_M_screen_y_q_4\ : std_logic;
signal \this_ppu.M_state_qZ0Z_6\ : std_logic;
signal \this_ppu.m68_0_a2_2_cascade_\ : std_logic;
signal \this_ppu.M_state_q_ns_7\ : std_logic;
signal \M_this_ppu_vga_is_drawing_cascade_\ : std_logic;
signal \this_ppu_M_screen_y_q_5\ : std_logic;
signal \this_ppu_M_screen_y_q_6\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c1\ : std_logic;
signal \M_this_scroll_qZ0Z_9\ : std_logic;
signal \M_this_scroll_qZ0Z_15\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_ac0_11\ : std_logic;
signal \M_this_scroll_qZ0Z_12\ : std_logic;
signal \this_ppu.un1_M_surface_x_q_c4\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_2\ : std_logic;
signal \M_this_map_ram_read_data_2\ : std_logic;
signal \M_this_ppu_spr_addr_8\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \this_ppu.M_screen_y_q_RNICCMV8Z0Z_0\ : std_logic;
signal \this_ppu.offset_y\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1\ : std_logic;
signal \this_ppu.M_surface_y_qZ0Z_1\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_0\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2\ : std_logic;
signal \this_ppu.M_surface_y_qZ0Z_2\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_1\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3\ : std_logic;
signal \M_this_ppu_map_addr_5\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_2\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4\ : std_logic;
signal \M_this_ppu_map_addr_6\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_3\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5\ : std_logic;
signal \M_this_ppu_map_addr_7\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_4\ : std_logic;
signal \this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6\ : std_logic;
signal \M_this_ppu_map_addr_8\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_5\ : std_logic;
signal \this_ppu.un1_M_surface_y_d_cry_6\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_7\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \M_this_ppu_map_addr_9\ : std_logic;
signal \M_this_ppu_vram_addr_7\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_1\ : std_logic;
signal \M_this_ppu_vga_is_drawing\ : std_logic;
signal \this_ppu.M_screen_y_qZ0Z_2\ : std_logic;
signal \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0\ : std_logic;
signal \M_this_oam_ram_read_data_12\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_12\ : std_logic;
signal \this_delay_clk.M_pipe_qZ0Z_3\ : std_logic;
signal \N_1256_0\ : std_logic;
signal \M_this_oam_ram_read_data_16\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_16\ : std_logic;
signal \M_this_oam_ram_read_data_17\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_17\ : std_logic;
signal \M_this_oam_ram_read_data_18\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_18\ : std_logic;
signal \M_this_oam_ram_read_data_27\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_27\ : std_logic;
signal \M_this_ctrl_flags_qZ0Z_6\ : std_logic;
signal \M_this_oam_ram_read_data_13\ : std_logic;
signal \this_ppu.M_state_qZ0Z_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_write_data_13\ : std_logic;
signal \M_this_oam_address_qZ0Z_1\ : std_logic;
signal \M_this_oam_address_qZ0Z_0\ : std_logic;
signal \N_222_0\ : std_logic;
signal \N_1248_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_2\ : std_logic;
signal \M_this_spr_ram_write_en_0_i_1_0_cascade_\ : std_logic;
signal \this_spr_ram.mem_WE_2\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lt8_0_cascade_\ : std_logic;
signal \this_ppu.offset_x\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_8\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_9\ : std_logic;
signal \this_ppu.M_surface_x_qZ0Z_1\ : std_logic;
signal \M_this_ppu_spr_addr_1\ : std_logic;
signal \this_ppu.offset_x_cry_0\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_10\ : std_logic;
signal \this_ppu.M_surface_x_qZ0Z_2\ : std_logic;
signal \M_this_ppu_spr_addr_2\ : std_logic;
signal \this_ppu.offset_x_cry_1\ : std_logic;
signal \M_this_ppu_map_addr_0\ : std_logic;
signal \this_ppu.offset_x_3\ : std_logic;
signal \this_ppu.offset_x_cry_2\ : std_logic;
signal \M_this_ppu_map_addr_1\ : std_logic;
signal \this_ppu.offset_x_4\ : std_logic;
signal \this_ppu.offset_x_cry_3\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_13\ : std_logic;
signal \M_this_ppu_map_addr_2\ : std_logic;
signal \this_ppu.offset_x_5\ : std_logic;
signal \this_ppu.offset_x_cry_4\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_14\ : std_logic;
signal \M_this_ppu_map_addr_3\ : std_logic;
signal \this_ppu.offset_x_6\ : std_logic;
signal \this_ppu.offset_x_cry_5\ : std_logic;
signal \M_this_ppu_map_addr_4\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_15\ : std_logic;
signal \this_ppu.offset_x_cry_6\ : std_logic;
signal \this_ppu.offset_x_7\ : std_logic;
signal \M_this_scroll_qZ0Z_0\ : std_logic;
signal \M_this_scroll_qZ0Z_1\ : std_logic;
signal \M_this_scroll_qZ0Z_2\ : std_logic;
signal \M_this_scroll_qZ0Z_3\ : std_logic;
signal \M_this_scroll_qZ0Z_4\ : std_logic;
signal \M_this_scroll_qZ0Z_5\ : std_logic;
signal \M_this_scroll_qZ0Z_6\ : std_logic;
signal \M_this_scroll_qZ0Z_7\ : std_logic;
signal \bfn_15_19_0_\ : std_logic;
signal \M_this_data_count_q_cry_0_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_0\ : std_logic;
signal \M_this_data_count_q_cry_1_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_1\ : std_logic;
signal \M_this_data_count_q_cry_2_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_2\ : std_logic;
signal \M_this_data_count_q_cry_3\ : std_logic;
signal \M_this_data_count_q_cry_4\ : std_logic;
signal \M_this_data_count_q_cry_5\ : std_logic;
signal \M_this_data_count_q_cry_6_THRU_CO\ : std_logic;
signal \M_this_data_count_q_cry_6\ : std_logic;
signal \M_this_data_count_q_cry_7\ : std_logic;
signal \bfn_15_20_0_\ : std_logic;
signal \M_this_data_count_q_cry_8\ : std_logic;
signal \M_this_data_count_q_cry_9\ : std_logic;
signal \M_this_data_count_q_cry_10\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \M_this_data_count_q_cry_11\ : std_logic;
signal \M_this_data_count_q_cry_12\ : std_logic;
signal port_enb_c : std_logic;
signal \M_this_delay_clk_out_0\ : std_logic;
signal \M_this_data_count_q_s_8\ : std_logic;
signal \N_92\ : std_logic;
signal \M_this_data_count_qZ0Z_8\ : std_logic;
signal \M_this_data_count_q_cry_3_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_4\ : std_logic;
signal \M_this_data_count_q_cry_4_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_5\ : std_logic;
signal \M_this_data_count_q_cry_8_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_9\ : std_logic;
signal \this_start_data_delay.M_last_qZ0\ : std_logic;
signal \N_685_i_cascade_\ : std_logic;
signal \M_this_data_count_qZ0Z_2\ : std_logic;
signal \M_this_data_count_qZ0Z_1\ : std_logic;
signal \M_this_data_count_qZ0Z_3\ : std_logic;
signal \M_this_data_count_qZ0Z_0\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_1\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_4\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_0\ : std_logic;
signal \M_this_map_ram_read_data_0\ : std_logic;
signal \M_this_ppu_spr_addr_6\ : std_logic;
signal \this_ppu.oam_cache.mem_0\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_1\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_2\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8\ : std_logic;
signal \this_vga_signals.M_vcounter_d7lto9_i_a2_1\ : std_logic;
signal port_nmib_1_i : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_11\ : std_logic;
signal \this_ppu.oam_cache.mem_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_11\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_12\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_i_12\ : std_logic;
signal \this_ppu.oam_cache.mem_8\ : std_logic;
signal \this_ppu.M_oam_cache_read_data_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_0\ : std_logic;
signal \this_vga_signals.N_3_1_cascade_\ : std_logic;
signal \this_vga_signals.g0_41_N_2L1\ : std_logic;
signal \this_vga_signals.g0_41_N_4L5_cascade_\ : std_logic;
signal \this_vga_signals.g0_41_1\ : std_logic;
signal \M_this_vga_ramdac_en\ : std_logic;
signal \this_vga_signals.mult1_un82_sum_c3_0_0_0_1\ : std_logic;
signal \M_this_vga_signals_address_7\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_\ : std_logic;
signal \this_vga_signals.N_17_i\ : std_logic;
signal \M_this_data_count_q_s_10\ : std_logic;
signal \M_this_data_count_q_cry_11_THRU_CO\ : std_logic;
signal \M_this_data_count_q_s_13\ : std_logic;
signal \M_this_data_count_q_cry_10_THRU_CO\ : std_logic;
signal \M_this_data_count_qZ0Z_7\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_12\ : std_logic;
signal \M_this_data_count_qZ0Z_11\ : std_logic;
signal \M_this_data_count_qZ0Z_13\ : std_logic;
signal \M_this_data_count_qZ0Z_10\ : std_logic;
signal \this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11\ : std_logic;
signal \M_this_data_count_q_cry_5_THRU_CO\ : std_logic;
signal \N_685_i\ : std_logic;
signal \M_this_data_count_qZ0Z_6\ : std_logic;
signal \M_this_ctrl_flags_qZ0Z_5\ : std_logic;
signal \M_this_ctrl_flags_qZ0Z_7\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_5\ : std_logic;
signal \M_this_spr_address_qZ0Z_0\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_spr_address_q_cry_0\ : std_logic;
signal \M_this_spr_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_spr_address_q_cry_1\ : std_logic;
signal \M_this_spr_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_spr_address_q_cry_2\ : std_logic;
signal \M_this_spr_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_spr_address_q_cry_3\ : std_logic;
signal \M_this_spr_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_spr_address_q_cry_4\ : std_logic;
signal \M_this_spr_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_5\ : std_logic;
signal \M_this_spr_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_spr_address_q_cry_6\ : std_logic;
signal \un1_M_this_spr_address_q_cry_7\ : std_logic;
signal \M_this_spr_address_qZ0Z_8\ : std_logic;
signal \bfn_17_13_0_\ : std_logic;
signal \M_this_spr_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_8\ : std_logic;
signal \M_this_spr_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_9\ : std_logic;
signal \un1_M_this_spr_address_q_cry_10\ : std_logic;
signal \un1_M_this_spr_address_q_cry_11\ : std_logic;
signal \un1_M_this_spr_address_q_cry_12\ : std_logic;
signal \M_this_spr_ram_write_en_0_i_1\ : std_logic;
signal \this_vga_signals.M_vcounter_d8\ : std_logic;
signal \this_vga_signals.M_hcounter_d7_0\ : std_logic;
signal \this_vga_signals.m43_5\ : std_logic;
signal this_vga_signals_vsync_1_i : std_logic;
signal \N_52_0\ : std_logic;
signal \N_58_0\ : std_logic;
signal \this_ppu.line_clk.M_last_qZ0\ : std_logic;
signal \this_vga_signals.GZ0Z_424\ : std_logic;
signal \this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9\ : std_logic;
signal \this_ppu.oam_cache.mem_1\ : std_logic;
signal \this_vga_signals.vvisibility_0_cascade_\ : std_logic;
signal \this_vga_signals.vvisibility\ : std_logic;
signal \this_vga_signals.g0_0_i_0_1\ : std_logic;
signal \this_vga_signals.N_10_i_cascade_\ : std_logic;
signal \this_vga_signals.g2_1_2\ : std_logic;
signal \this_vga_signals.N_10_i_0\ : std_logic;
signal \this_vga_signals.g0_0_i_0_cascade_\ : std_logic;
signal \this_vga_signals.if_m5_i_0_0\ : std_logic;
signal \this_vga_signals.mult1_un68_sum_c3_0_0_0\ : std_logic;
signal \this_vga_signals.if_N_10_0_0_0\ : std_logic;
signal \this_vga_signals.g0_1_0_3\ : std_logic;
signal \this_vga_signals.g0_1_1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\ : std_logic;
signal \this_vga_signals.g0_41_N_3L3_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_x0_cascade_\ : std_logic;
signal \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_\ : std_logic;
signal \this_vga_signals.g0_41_N_4L5_1\ : std_logic;
signal \N_6_i\ : std_logic;
signal \this_vga_signals.g0_1_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c2_0_0\ : std_logic;
signal \this_vga_signals.g1_4\ : std_logic;
signal \this_vga_signals.g1_0_0_0\ : std_logic;
signal \this_vga_signals.g1_0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.N_10\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_2_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_\ : std_logic;
signal \this_vga_signals.N_5_i_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_i_x2_1\ : std_logic;
signal \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\ : std_logic;
signal \this_spr_ram.mem_WE_8\ : std_logic;
signal \this_vga_signals.m43_4\ : std_logic;
signal \this_vga_signals.vaddress_c3_d_0\ : std_logic;
signal \this_vga_signals.g0_1_0_1\ : std_logic;
signal \this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_\ : std_logic;
signal \this_vga_signals.CO0_0_i_i_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_c5_a0_0_cascade_\ : std_logic;
signal \this_vga_signals.vaddress_9_cascade_\ : std_logic;
signal \this_vga_signals.g1_3_0_cascade_\ : std_logic;
signal \this_vga_signals.N_5_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_c3_0_0_0\ : std_logic;
signal \this_vga_signals.N_4_1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c3_x1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0_cascade_\ : std_logic;
signal \this_vga_signals.g1_1_0_0_cascade_\ : std_logic;
signal \this_vga_signals.N_20_0\ : std_logic;
signal \this_vga_signals.g0_2_0_3_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_0_1_0\ : std_logic;
signal \this_vga_signals.g0_0_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4\ : std_logic;
signal \this_vga_signals.g0_2_0_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_4\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0\ : std_logic;
signal \this_vga_signals.g0_6_0\ : std_logic;
signal \this_vga_signals.g0_0_0_1\ : std_logic;
signal \this_vga_signals.g0_5_5_N_2L1\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0 : std_logic;
signal \this_vga_signals.g0_5_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3\ : std_logic;
signal \this_vga_signals.g1_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_d_0\ : std_logic;
signal \this_vga_signals.g0_1_0_cascade_\ : std_logic;
signal \this_vga_signals.N_7_1_0_2\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\ : std_logic;
signal \this_vga_signals.g3_1\ : std_logic;
signal \this_vga_signals.g1_3\ : std_logic;
signal \this_vga_signals.N_7_1_0_0\ : std_logic;
signal \this_vga_signals.g0_1_0_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_ns\ : std_logic;
signal \this_vga_signals.g1_0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_c2_0\ : std_logic;
signal \this_vga_signals.g0_29_1\ : std_logic;
signal \this_vga_signals.g1_0_cascade_\ : std_logic;
signal this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0 : std_logic;
signal \this_vga_signals.g0_3\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_6\ : std_logic;
signal \M_this_reset_cond_out_0\ : std_logic;
signal rst_n_c : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_7\ : std_logic;
signal \this_reset_cond.M_stage_qZ0Z_8\ : std_logic;
signal \this_spr_ram.mem_WE_10\ : std_logic;
signal \this_vga_signals.N_12_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_4\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_5\ : std_logic;
signal \this_vga_signals.vaddress_c2_cascade_\ : std_logic;
signal \this_vga_signals.N_7_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0\ : std_logic;
signal \this_vga_signals.g0_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_x0\ : std_logic;
signal \this_vga_signals.vaddress_ac0_9_0_a0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_\ : std_logic;
signal \this_vga_signals.g0_5_5\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_3\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_2\ : std_logic;
signal \this_vga_signals.N_5_i_1\ : std_logic;
signal \this_vga_signals.N_5786_0_0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x0\ : std_logic;
signal \this_vga_signals.mult1_un47_sum_axbxc3_x1\ : std_logic;
signal \this_vga_signals.CO0_0_i_i\ : std_logic;
signal \this_vga_signals.N_12_0\ : std_logic;
signal \this_vga_signals.N_12_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_axb1_0_1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_x0\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_ns\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axbxc3_1\ : std_logic;
signal \this_vga_signals.g0_2_0_1\ : std_logic;
signal \this_vga_signals.mult1_un54_sum_axb1_out_0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\ : std_logic;
signal port_rw_in : std_logic;
signal \M_this_state_d_0_sqmuxa_2_cascade_\ : std_logic;
signal \this_start_data_delay.N_233_0_cascade_\ : std_logic;
signal \N_164\ : std_logic;
signal \this_vga_signals.g1_3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6\ : std_logic;
signal \this_spr_ram.mem_WE_6\ : std_logic;
signal \M_this_spr_address_qZ0Z_12\ : std_logic;
signal \M_this_spr_address_qZ0Z_11\ : std_logic;
signal \M_this_spr_address_qZ0Z_13\ : std_logic;
signal \M_this_spr_ram_write_en_0_i_1_0\ : std_logic;
signal \this_spr_ram.mem_WE_4\ : std_logic;
signal \M_this_spr_ram_write_data_3\ : std_logic;
signal \this_ppu.oam_cache.M_oam_cache_read_data_1\ : std_logic;
signal \M_this_map_ram_read_data_1\ : std_logic;
signal \this_ppu.M_state_q_inv_1\ : std_logic;
signal \M_this_ppu_spr_addr_7\ : std_logic;
signal \M_this_spr_ram_write_data_1\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_c3_0\ : std_logic;
signal \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_\ : std_logic;
signal \this_vga_signals.N_14\ : std_logic;
signal \this_vga_signals.g1_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_5\ : std_logic;
signal \this_vga_signals.N_7_1_0_3_cascade_\ : std_logic;
signal \this_vga_signals.G_5_i_o2_0_1\ : std_logic;
signal \this_vga_signals.vaddress_8\ : std_logic;
signal \this_vga_signals.vaddress_9\ : std_logic;
signal \this_vga_signals.N_19_0_0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_6\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_9\ : std_logic;
signal \this_vga_signals.m47_0_0\ : std_logic;
signal \this_vga_signals.m47_0_1_cascade_\ : std_logic;
signal \this_vga_signals_M_vcounter_q_6\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_4\ : std_logic;
signal \this_vga_signals.SUM_2_cascade_\ : std_logic;
signal \this_vga_signals.g0_0_i_a7_1\ : std_logic;
signal \N_88\ : std_logic;
signal port_address_in_5 : std_logic;
signal port_address_in_7 : std_logic;
signal port_address_in_3 : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\ : std_logic;
signal \this_vga_signals.M_vcounter_q_4_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_5_repZ0Z1\ : std_logic;
signal \this_vga_signals.vaddress_7\ : std_logic;
signal \this_vga_signals.vaddress_6\ : std_logic;
signal \this_vga_signals.vaddress_5\ : std_logic;
signal \this_vga_signals.vaddress_7_cascade_\ : std_logic;
signal \this_vga_signals.SUM_2\ : std_logic;
signal \this_vga_signals.if_m2_0\ : std_logic;
signal \this_start_data_delay.N_345_cascade_\ : std_logic;
signal \this_start_data_delay.N_284_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_\ : std_logic;
signal \this_start_data_delay.N_23_1_0_cascade_\ : std_logic;
signal \this_start_data_delay.N_339_cascade_\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6\ : std_logic;
signal \M_this_substate_qZ0\ : std_logic;
signal \this_start_data_delay.N_467\ : std_logic;
signal \this_start_data_delay.N_386_cascade_\ : std_logic;
signal port_address_in_1 : std_logic;
signal \this_start_data_delay.N_380\ : std_logic;
signal \this_start_data_delay.N_341\ : std_logic;
signal \M_this_spr_ram_write_data_2\ : std_logic;
signal \dma_axb0_cascade_\ : std_logic;
signal dma_0 : std_logic;
signal dma_axb3 : std_logic;
signal \this_vga_signals.vaddress_c2\ : std_logic;
signal \this_vga_signals.N_13\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_7\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\ : std_logic;
signal \this_vga_signals_M_vcounter_q_8\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\ : std_logic;
signal \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\ : std_logic;
signal \this_vga_signals.N_933_0\ : std_logic;
signal \this_vga_signals.N_1188_g\ : std_logic;
signal \N_422_2_cascade_\ : std_logic;
signal \N_458_i\ : std_logic;
signal \this_vga_signals.M_vcounter_q_6_repZ0Z1\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_8\ : std_logic;
signal \this_vga_signals.M_vcounter_qZ0Z_9\ : std_logic;
signal \this_vga_signals.M_vcounter_q_fastZ0Z_7\ : std_logic;
signal \this_vga_signals.mult1_un40_sum_ac0_3_1_1\ : std_logic;
signal \this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3\ : std_logic;
signal \this_start_data_delay.N_424\ : std_logic;
signal \M_this_spr_ram_write_data_0\ : std_logic;
signal \M_this_state_qZ0Z_11\ : std_logic;
signal \this_start_data_delay.N_245_0_cascade_\ : std_logic;
signal un20_i_a4_0_a2_0_a2_1 : std_logic;
signal \M_this_state_qZ0Z_13\ : std_logic;
signal un20_i_a4_0_a2_2 : std_logic;
signal \N_241_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_\ : std_logic;
signal \this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0\ : std_logic;
signal \M_this_state_qZ0Z_12\ : std_logic;
signal \this_start_data_delay.N_245_0\ : std_logic;
signal \M_this_state_qZ0Z_7\ : std_logic;
signal \M_this_state_qZ0Z_8\ : std_logic;
signal port_address_in_2 : std_logic;
signal port_address_in_6 : std_logic;
signal \this_vga_signals_M_this_state_d28_0_a2_0_1\ : std_logic;
signal \N_1264_0\ : std_logic;
signal \this_start_data_delay.N_387\ : std_logic;
signal port_address_in_0 : std_logic;
signal port_address_in_4 : std_logic;
signal \this_start_data_delay.N_337_cascade_\ : std_logic;
signal \this_start_data_delay.N_386\ : std_logic;
signal \M_this_state_qZ0Z_6\ : std_logic;
signal \M_this_state_qZ0Z_5\ : std_logic;
signal \this_start_data_delay.N_239_0\ : std_logic;
signal \M_this_state_qZ0Z_3\ : std_logic;
signal \M_this_state_qZ0Z_2\ : std_logic;
signal \M_this_state_qZ0Z_1\ : std_logic;
signal \this_start_data_delay.N_420_3\ : std_logic;
signal \this_start_data_delay.N_23_1_0\ : std_logic;
signal \this_start_data_delay.N_344_cascade_\ : std_logic;
signal \N_465\ : std_logic;
signal \this_start_data_delay.N_246_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0\ : std_logic;
signal \M_last_q_RNIE8SF1\ : std_logic;
signal \M_this_ext_address_qZ0Z_0\ : std_logic;
signal \bfn_21_24_0_\ : std_logic;
signal \M_this_ext_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_ext_address_q_cry_0\ : std_logic;
signal \M_this_ext_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_ext_address_q_cry_1\ : std_logic;
signal \M_this_ext_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_ext_address_q_cry_2\ : std_logic;
signal \M_this_ext_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_ext_address_q_cry_3\ : std_logic;
signal \M_this_ext_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_ext_address_q_cry_4\ : std_logic;
signal \M_this_ext_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_ext_address_q_cry_5\ : std_logic;
signal \M_this_ext_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_ext_address_q_cry_6\ : std_logic;
signal \un1_M_this_ext_address_q_cry_7\ : std_logic;
signal \M_this_ext_address_qZ0Z_8\ : std_logic;
signal \bfn_21_25_0_\ : std_logic;
signal \M_this_ext_address_qZ0Z_9\ : std_logic;
signal \un1_M_this_ext_address_q_cry_8\ : std_logic;
signal \M_this_ext_address_qZ0Z_10\ : std_logic;
signal \un1_M_this_ext_address_q_cry_9\ : std_logic;
signal \M_this_ext_address_qZ0Z_11\ : std_logic;
signal \un1_M_this_ext_address_q_cry_10\ : std_logic;
signal \M_this_ext_address_qZ0Z_12\ : std_logic;
signal \un1_M_this_ext_address_q_cry_11\ : std_logic;
signal \M_this_ext_address_qZ0Z_13\ : std_logic;
signal \un1_M_this_ext_address_q_cry_12\ : std_logic;
signal \M_this_ext_address_qZ0Z_14\ : std_logic;
signal \un1_M_this_ext_address_q_cry_13\ : std_logic;
signal \N_295\ : std_logic;
signal \un1_M_this_ext_address_q_cry_14\ : std_logic;
signal \M_this_ext_address_qZ0Z_15\ : std_logic;
signal \this_start_data_delay.N_231_0\ : std_logic;
signal \M_this_reset_cond_out_g_0\ : std_logic;
signal \this_start_data_delay.N_227_0\ : std_logic;
signal \this_start_data_delay.N_242_0\ : std_logic;
signal \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_\ : std_logic;
signal \N_220_0\ : std_logic;
signal \M_this_state_qZ0Z_10\ : std_logic;
signal \N_930\ : std_logic;
signal \M_this_state_qZ0Z_9\ : std_logic;
signal \M_this_state_qZ0Z_4\ : std_logic;
signal \this_start_data_delay.N_332\ : std_logic;
signal port_data_c_0 : std_logic;
signal \M_this_map_ram_write_data_0\ : std_logic;
signal led_c_1 : std_logic;
signal \N_466\ : std_logic;
signal led_c_7 : std_logic;
signal port_data_c_3 : std_logic;
signal \M_this_map_ram_write_data_3\ : std_logic;
signal port_data_c_1 : std_logic;
signal \M_this_map_ram_write_data_1\ : std_logic;
signal port_data_c_2 : std_logic;
signal \M_this_map_ram_write_data_2\ : std_logic;
signal port_data_c_4 : std_logic;
signal \M_this_map_ram_write_data_4\ : std_logic;
signal port_data_c_6 : std_logic;
signal \M_this_map_ram_write_data_6\ : std_logic;
signal port_data_c_5 : std_logic;
signal \M_this_map_ram_write_data_5\ : std_logic;
signal port_data_c_7 : std_logic;
signal \M_this_map_ram_write_data_7\ : std_logic;
signal \M_this_state_d_0_sqmuxa\ : std_logic;
signal \M_this_map_address_qZ0Z_0\ : std_logic;
signal \bfn_26_25_0_\ : std_logic;
signal \M_this_map_address_qZ0Z_1\ : std_logic;
signal \un1_M_this_map_address_q_cry_0\ : std_logic;
signal \M_this_map_address_qZ0Z_2\ : std_logic;
signal \un1_M_this_map_address_q_cry_1\ : std_logic;
signal \M_this_map_address_qZ0Z_3\ : std_logic;
signal \un1_M_this_map_address_q_cry_2\ : std_logic;
signal \M_this_map_address_qZ0Z_4\ : std_logic;
signal \un1_M_this_map_address_q_cry_3\ : std_logic;
signal \M_this_map_address_qZ0Z_5\ : std_logic;
signal \un1_M_this_map_address_q_cry_4\ : std_logic;
signal \M_this_map_address_qZ0Z_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_5\ : std_logic;
signal \M_this_map_address_qZ0Z_7\ : std_logic;
signal \un1_M_this_map_address_q_cry_6\ : std_logic;
signal \un1_M_this_map_address_q_cry_7\ : std_logic;
signal \M_this_map_address_qZ0Z_8\ : std_logic;
signal \bfn_26_26_0_\ : std_logic;
signal \N_93\ : std_logic;
signal \un1_M_this_map_address_q_cry_8\ : std_logic;
signal \M_this_map_address_qZ0Z_9\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_0_c_g : std_logic;
signal \N_527_g\ : std_logic;

signal clk_wire : std_logic;
signal debug_wire : std_logic_vector(1 downto 0);
signal hblank_wire : std_logic;
signal hsync_wire : std_logic;
signal led_wire : std_logic_vector(7 downto 0);
signal port_clk_wire : std_logic;
signal port_data_wire : std_logic_vector(7 downto 0);
signal port_data_rw_wire : std_logic;
signal port_dmab_wire : std_logic;
signal port_enb_wire : std_logic;
signal port_nmib_wire : std_logic;
signal rgb_wire : std_logic_vector(5 downto 0);
signal rst_n_wire : std_logic;
signal vblank_wire : std_logic;
signal vsync_wire : std_logic;
signal \this_map_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \this_vram.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \this_vram.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    clk_wire <= clk;
    debug <= debug_wire;
    hblank <= hblank_wire;
    hsync <= hsync_wire;
    led <= led_wire;
    port_clk_wire <= port_clk;
    port_data_wire <= port_data;
    port_data_rw <= port_data_rw_wire;
    port_dmab <= port_dmab_wire;
    port_enb_wire <= port_enb;
    port_nmib <= port_nmib_wire;
    rgb <= rgb_wire;
    rst_n_wire <= rst_n;
    vblank <= vblank_wire;
    vsync <= vsync_wire;
    \M_this_map_ram_read_data_3\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_2\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_1\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_0\ <= \this_map_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&\N__23300\&\N__22445\&\N__22505\&\N__22556\&\N__22613\&\N__25064\&\N__24110\&\N__24188\&\N__24266\&\N__24329\;
    \this_map_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&\N__39461\&\N__39560\&\N__39590\&\N__39617\&\N__38375\&\N__38405\&\N__38432\&\N__38462\&\N__38492\&\N__38519\;
    \this_map_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&\N__37772\&'0'&'0'&'0'&\N__37535\&'0'&'0'&'0'&\N__37658\&'0'&'0'&'0'&\N__38024\&'0';
    \M_this_map_ram_read_data_7\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_map_ram_read_data_6\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_map_ram_read_data_5\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_map_ram_read_data_4\ <= \this_map_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_map_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&\N__23293\&\N__22439\&\N__22499\&\N__22546\&\N__22607\&\N__25058\&\N__24104\&\N__24182\&\N__24260\&\N__24319\;
    \this_map_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&\N__39455\&\N__39554\&\N__39584\&\N__39611\&\N__38369\&\N__38399\&\N__38426\&\N__38456\&\N__38486\&\N__38513\;
    \this_map_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_map_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&\N__38636\&'0'&'0'&'0'&\N__37259\&'0'&'0'&'0'&\N__38780\&'0'&'0'&'0'&\N__37406\&'0';
    \M_this_oam_ram_read_data_15\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_14\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_13\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_12\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_11\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_10\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_9\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_8\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_7\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_6\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_5\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_4\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_3\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_2\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_1\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_0\ <= \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__18947\&\N__18680\&\N__18260\&\N__18349\&\N__18425\&\N__18551\;
    \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__17198\&\N__17231\&\N__19520\&\N__19481\&\N__19604\&\N__19568\;
    \this_oam_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\ <= \N__15080\&\N__14846\&\N__15086\&\N__16637\&\N__17549\&\N__16649\&\N__17576\&\N__15038\&\N__15206\&\N__14978\&\N__15212\&\N__17567\&\N__15023\&\N__17594\&\N__17627\&\N__19229\;
    \M_this_oam_ram_read_data_31\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(15);
    \M_this_oam_ram_read_data_30\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(14);
    \M_this_oam_ram_read_data_29\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(13);
    \M_this_oam_ram_read_data_28\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(12);
    \M_this_oam_ram_read_data_27\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \M_this_oam_ram_read_data_26\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(10);
    \M_this_oam_ram_read_data_25\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(9);
    \M_this_oam_ram_read_data_24\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(8);
    \M_this_oam_ram_read_data_23\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(7);
    \M_this_oam_ram_read_data_22\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(6);
    \M_this_oam_ram_read_data_21\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(5);
    \M_this_oam_ram_read_data_20\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(4);
    \M_this_oam_ram_read_data_19\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \M_this_oam_ram_read_data_18\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(2);
    \M_this_oam_ram_read_data_17\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(1);
    \M_this_oam_ram_read_data_16\ <= \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__18941\&\N__18674\&\N__18254\&\N__18336\&\N__18419\&\N__18545\;
    \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__17192\&\N__17225\&\N__19514\&\N__19475\&\N__19598\&\N__19562\;
    \this_oam_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\ <= \N__16601\&\N__15464\&\N__15452\&\N__17756\&\N__15470\&\N__19406\&\N__17747\&\N__15446\&\N__16790\&\N__15149\&\N__16802\&\N__17606\&\N__17768\&\N__15074\&\N__15458\&\N__15158\;
    \this_ppu.oam_cache.mem_15\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(15);
    \this_ppu.oam_cache.mem_14\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(14);
    \this_ppu.oam_cache.mem_13\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(13);
    \this_ppu.oam_cache.mem_12\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(12);
    \this_ppu.oam_cache.mem_11\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_ppu.oam_cache.mem_10\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(10);
    \this_ppu.oam_cache.mem_9\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(9);
    \this_ppu.oam_cache.mem_8\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(8);
    \this_ppu.oam_cache.mem_7\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(7);
    \this_ppu.oam_cache.mem_6\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(6);
    \this_ppu.oam_cache.mem_5\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(5);
    \this_ppu.oam_cache.mem_4\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(4);
    \this_ppu.oam_cache.mem_3\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_ppu.oam_cache.mem_2\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_1\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_0\ <= \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18185\&\N__14735\&\N__14720\&\N__14699\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__13709\&\N__13412\&\N__13367\&\N__13454\;
    \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\ <= \N__13295\&\N__13319\&\N__23783\&\N__23009\&\N__19181\&\N__13220\&\N__13238\&\N__13259\&\N__13631\&\N__13283\&\N__13655\&\N__13643\&\N__13289\&\N__13667\&\N__13619\&\N__13673\;
    \this_ppu.oam_cache.mem_18\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(2);
    \this_ppu.oam_cache.mem_17\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(1);
    \this_ppu.oam_cache.mem_16\ <= \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\(0);
    \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__18179\&\N__14729\&\N__14714\&\N__14693\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__13701\&\N__13404\&\N__13361\&\N__13446\;
    \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\ <= \N__15053\&\N__14831\&\N__15170\&\N__15191\&\N__23336\&\N__14855\&\N__14876\&\N__14903\&\N__14927\&\N__14750\&\N__14756\&\N__15101\&\N__15140\&\N__23369\&\N__23417\&\N__23459\;
    \this_spr_ram.mem_out_bus0_1\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_0\ <= \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\ <= \N__20314\&\N__20580\&\N__22983\&\N__32561\&\N__26290\&\N__15846\&\N__16008\&\N__17429\&\N__24483\&\N__24797\&\N__20147\;
    \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\ <= \N__28912\&\N__29101\&\N__29349\&\N__29570\&\N__27113\&\N__27334\&\N__27521\&\N__27806\&\N__28049\&\N__28207\&\N__28414\;
    \this_spr_ram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32373\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35085\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus0_3\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus0_2\ <= \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\ <= \N__20315\&\N__20581\&\N__22921\&\N__32535\&\N__26219\&\N__15827\&\N__16065\&\N__17455\&\N__24506\&\N__24738\&\N__20148\;
    \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\ <= \N__28903\&\N__29100\&\N__29348\&\N__29569\&\N__27073\&\N__27280\&\N__27550\&\N__27802\&\N__28055\&\N__28236\&\N__28477\;
    \this_spr_ram.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32818\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34276\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_1\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_0\ <= \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\ <= \N__20350\&\N__20619\&\N__22993\&\N__32562\&\N__26289\&\N__15872\&\N__16088\&\N__17475\&\N__24501\&\N__24814\&\N__20176\;
    \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\ <= \N__28902\&\N__29121\&\N__29354\&\N__29576\&\N__27130\&\N__27281\&\N__27497\&\N__27795\&\N__28048\&\N__28257\&\N__28495\;
    \this_spr_ram.mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32374\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35097\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus1_3\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus1_2\ <= \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\ <= \N__20351\&\N__20620\&\N__22987\&\N__32563\&\N__26294\&\N__15873\&\N__16089\&\N__17489\&\N__24525\&\N__24801\&\N__20177\;
    \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\ <= \N__28877\&\N__29028\&\N__29353\&\N__29575\&\N__27137\&\N__27282\&\N__27525\&\N__27775\&\N__28006\&\N__28269\&\N__28506\;
    \this_spr_ram.mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32819\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34282\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_1\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_0\ <= \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\ <= \N__20405\&\N__20648\&\N__22994\&\N__32588\&\N__26263\&\N__15888\&\N__16109\&\N__17501\&\N__24536\&\N__24836\&\N__20146\;
    \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\ <= \N__28868\&\N__29047\&\N__29286\&\N__29571\&\N__27134\&\N__27316\&\N__27566\&\N__27742\&\N__28005\&\N__28274\&\N__28505\;
    \this_spr_ram.mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32396\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35102\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus2_3\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus2_2\ <= \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\ <= \N__20401\&\N__20647\&\N__22989\&\N__32587\&\N__26300\&\N__15887\&\N__16108\&\N__17497\&\N__24502\&\N__24832\&\N__20145\;
    \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\ <= \N__28869\&\N__29080\&\N__29341\&\N__29546\&\N__27120\&\N__27317\&\N__27496\&\N__27744\&\N__28050\&\N__28270\&\N__28491\;
    \this_spr_ram.mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32814\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34277\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_1\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_0\ <= \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\ <= \N__20393\&\N__20640\&\N__22988\&\N__32580\&\N__26220\&\N__15856\&\N__16101\&\N__17490\&\N__24548\&\N__24739\&\N__20198\;
    \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\ <= \N__28870\&\N__29081\&\N__29340\&\N__29550\&\N__27066\&\N__27319\&\N__27562\&\N__27743\&\N__28051\&\N__28262\&\N__28470\;
    \this_spr_ram.mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32392\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35098\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus3_3\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus3_2\ <= \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\ <= \N__20379\&\N__20627\&\N__22972\&\N__32579\&\N__26295\&\N__15854\&\N__16046\&\N__17479\&\N__24544\&\N__24825\&\N__20192\;
    \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\ <= \N__28900\&\N__29105\&\N__29311\&\N__29514\&\N__27106\&\N__27318\&\N__27555\&\N__27784\&\N__28031\&\N__28247\&\N__28469\;
    \this_spr_ram.mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32801\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34263\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_1\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_0\ <= \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\ <= \N__20359\&\N__20622\&\N__22971\&\N__32565\&\N__26296\&\N__15853\&\N__16091\&\N__17428\&\N__24537\&\N__24815\&\N__20178\;
    \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\ <= \N__28901\&\N__29122\&\N__29318\&\N__29515\&\N__27079\&\N__27343\&\N__27540\&\N__27785\&\N__28004\&\N__28223\&\N__28437\;
    \this_spr_ram.mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32385\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35089\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus4_3\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus4_2\ <= \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\ <= \N__20322\&\N__20588\&\N__22941\&\N__32564\&\N__26276\&\N__15893\&\N__16090\&\N__17463\&\N__24526\&\N__24802\&\N__20119\;
    \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\ <= \N__28911\&\N__29135\&\N__29285\&\N__29448\&\N__27033\&\N__27344\&\N__27463\&\N__27770\&\N__28037\&\N__28125\&\N__28429\;
    \this_spr_ram.mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32815\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34245\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_1\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_0\ <= \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\ <= \N__20352\&\N__20621\&\N__22940\&\N__32537\&\N__26279\&\N__15889\&\N__16073\&\N__17462\&\N__24510\&\N__24784\&\N__20155\;
    \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\ <= \N__28898\&\N__29142\&\N__29287\&\N__29572\&\N__27074\&\N__27336\&\N__27533\&\N__27771\&\N__28036\&\N__28191\&\N__28430\;
    \this_spr_ram.mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32375\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35072\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus5_3\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus5_2\ <= \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\ <= \N__20377\&\N__20623\&\N__22900\&\N__32536\&\N__26277\&\N__15880\&\N__16072\&\N__17443\&\N__24462\&\N__24758\&\N__20165\;
    \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\ <= \N__28899\&\N__29143\&\N__29288\&\N__29555\&\N__27075\&\N__27335\&\N__27553\&\N__27763\&\N__28032\&\N__28203\&\N__28465\;
    \this_spr_ram.mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32775\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34244\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_1\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_0\ <= \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\ <= \N__20378\&\N__20639\&\N__22859\&\N__32555\&\N__26278\&\N__15837\&\N__16047\&\N__17439\&\N__24443\&\N__24694\&\N__20185\;
    \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\ <= \N__28894\&\N__29147\&\N__29289\&\N__29551\&\N__27105\&\N__27320\&\N__27554\&\N__27762\&\N__28052\&\N__28235\&\N__28490\;
    \this_spr_ram.mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32360\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35051\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus6_3\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus6_2\ <= \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\ <= \N__20343\&\N__20612\&\N__22957\&\N__32556\&\N__26298\&\N__15822\&\N__15975\&\N__17350\&\N__24480\&\N__24770\&\N__20169\;
    \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\ <= \N__28890\&\N__29099\&\N__29350\&\N__29562\&\N__27083\&\N__27276\&\N__27551\&\N__27774\&\N__28041\&\N__28184\&\N__28459\;
    \this_spr_ram.mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32816\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34278\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_1\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_0\ <= \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\ <= \N__20389\&\N__20637\&\N__22967\&\N__32557\&\N__26299\&\N__15826\&\N__16006\&\N__17351\&\N__24481\&\N__24780\&\N__20196\;
    \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\ <= \N__28913\&\N__29098\&\N__29351\&\N__29573\&\N__27135\&\N__27333\&\N__27552\&\N__27772\&\N__28054\&\N__28243\&\N__28507\;
    \this_spr_ram.mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32372\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__35096\&'0'&'0'&'0';
    \this_spr_ram.mem_out_bus7_3\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(11);
    \this_spr_ram.mem_out_bus7_2\ <= \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\(3);
    \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\ <= \N__20400\&\N__20638\&\N__22982\&\N__32578\&\N__26297\&\N__15855\&\N__16007\&\N__17374\&\N__24482\&\N__24796\&\N__20197\;
    \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\ <= \N__28907\&\N__29120\&\N__29352\&\N__29574\&\N__27136\&\N__27312\&\N__27532\&\N__27773\&\N__28053\&\N__28261\&\N__28508\;
    \this_spr_ram.mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__32817\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__34283\&'0'&'0'&'0';
    \M_this_vram_read_data_3\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(3);
    \M_this_vram_read_data_2\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(2);
    \M_this_vram_read_data_1\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(1);
    \M_this_vram_read_data_0\ <= \this_vram.mem_mem_0_0_physical_RDATA_wire\(0);
    \this_vram.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&\N__26426\&\N__12728\&\N__13154\&\N__13127\&\N__13169\&\N__13019\&\N__12839\&\N__12983\;
    \this_vram.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&\N__23264\&\N__17003\&\N__17027\&\N__16844\&\N__17897\&\N__16904\&\N__16976\&\N__16946\;
    \this_vram.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \this_vram.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__17786\&\N__18692\&\N__17846\&\N__16694\;

    \this_map_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39418\,
            RE => \N__25718\,
            WCLKE => \N__38630\,
            WCLK => \N__39419\,
            WE => \N__25720\
        );

    \this_map_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_map_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_map_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_map_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_map_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_map_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39428\,
            RE => \N__25719\,
            WCLKE => \N__38625\,
            WCLK => \N__39429\,
            WE => \N__25721\
        );

    \this_oam_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39431\,
            RE => \N__25678\,
            WCLKE => \N__19391\,
            WCLK => \N__39432\,
            WE => \N__25680\
        );

    \this_oam_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_oam_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_oam_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_oam_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_oam_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_oam_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39433\,
            RE => \N__25679\,
            WCLKE => \N__19390\,
            WCLK => \N__39434\,
            WE => \N__25681\
        );

    \this_ppu.oam_cache.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39387\,
            RE => \N__25503\,
            WCLKE => \N__23950\,
            WCLK => \N__39388\,
            WE => \N__25599\
        );

    \this_ppu.oam_cache.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_ppu.oam_cache.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_ppu.oam_cache.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_ppu.oam_cache.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39400\,
            RE => \N__25543\,
            WCLKE => \N__24005\,
            WCLK => \N__39401\,
            WE => \N__25581\
        );

    \this_spr_ram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39298\,
            RE => \N__25722\,
            WCLKE => \N__16753\,
            WCLK => \N__39299\,
            WE => \N__25724\
        );

    \this_spr_ram.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39291\,
            RE => \N__25723\,
            WCLKE => \N__16757\,
            WCLK => \N__39292\,
            WE => \N__25766\
        );

    \this_spr_ram.mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39284\,
            RE => \N__25795\,
            WCLKE => \N__16774\,
            WCLK => \N__39285\,
            WE => \N__25580\
        );

    \this_spr_ram.mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_1_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_1_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39280\,
            RE => \N__25796\,
            WCLKE => \N__16778\,
            WCLK => \N__39281\,
            WE => \N__25797\
        );

    \this_spr_ram.mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39282\,
            RE => \N__25800\,
            WCLKE => \N__30722\,
            WCLK => \N__39283\,
            WE => \N__25799\
        );

    \this_spr_ram.mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_2_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_2_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39286\,
            RE => \N__25801\,
            WCLKE => \N__30718\,
            WCLK => \N__39287\,
            WE => \N__25798\
        );

    \this_spr_ram.mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39294\,
            RE => \N__25777\,
            WCLKE => \N__30113\,
            WCLK => \N__39295\,
            WE => \N__25788\
        );

    \this_spr_ram.mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_3_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_3_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39303\,
            RE => \N__25776\,
            WCLKE => \N__30109\,
            WCLK => \N__39304\,
            WE => \N__25787\
        );

    \this_spr_ram.mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39315\,
            RE => \N__25737\,
            WCLKE => \N__32246\,
            WCLK => \N__39314\,
            WE => \N__25765\
        );

    \this_spr_ram.mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_4_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_4_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39328\,
            RE => \N__25736\,
            WCLKE => \N__32245\,
            WCLK => \N__39329\,
            WE => \N__25764\
        );

    \this_spr_ram.mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39347\,
            RE => \N__25683\,
            WCLKE => \N__31837\,
            WCLK => \N__39348\,
            WE => \N__25684\
        );

    \this_spr_ram.mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_5_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_5_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39364\,
            RE => \N__25685\,
            WCLKE => \N__31838\,
            WCLK => \N__39365\,
            WE => \N__25717\
        );

    \this_spr_ram.mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39379\,
            RE => \N__25618\,
            WCLKE => \N__23557\,
            WCLK => \N__39380\,
            WE => \N__25625\
        );

    \this_spr_ram.mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_6_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_6_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39406\,
            RE => \N__25544\,
            WCLKE => \N__23564\,
            WCLK => \N__39407\,
            WE => \N__25582\
        );

    \this_spr_ram.mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_0_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_0_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39415\,
            RE => \N__25660\,
            WCLKE => \N__16714\,
            WCLK => \N__39416\,
            WE => \N__25601\
        );

    \this_spr_ram.mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_spr_ram.mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \this_spr_ram.mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \this_spr_ram.mem_mem_7_1_physical_WADDR_wire\,
            MASK => \this_spr_ram.mem_mem_7_1_physical_MASK_wire\,
            WDATA => \this_spr_ram.mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39425\,
            RE => \N__25661\,
            WCLKE => \N__16721\,
            WCLK => \N__39426\,
            WE => \N__25602\
        );

    \this_vram.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \this_vram.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \this_vram.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \this_vram.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \this_vram.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \this_vram.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__39372\,
            RE => \N__25515\,
            WCLKE => \N__20930\,
            WCLK => \N__39373\,
            WE => \N__25600\
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__40095\,
            GLOBALBUFFEROUTPUT => clk_0_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40097\,
            DIN => \N__40096\,
            DOUT => \N__40095\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__40097\,
            PADOUT => \N__40096\,
            PADIN => \N__40095\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40086\,
            DIN => \N__40085\,
            DOUT => \N__40084\,
            PACKAGEPIN => debug_wire(0)
        );

    \debug_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40086\,
            PADOUT => \N__40085\,
            PADIN => \N__40084\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \debug_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40077\,
            DIN => \N__40076\,
            DOUT => \N__40075\,
            PACKAGEPIN => debug_wire(1)
        );

    \debug_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40077\,
            PADOUT => \N__40076\,
            PADIN => \N__40075\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40068\,
            DIN => \N__40067\,
            DOUT => \N__40066\,
            PACKAGEPIN => hblank_wire
        );

    \hblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40068\,
            PADOUT => \N__40067\,
            PADIN => \N__40066\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12920\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \hsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40059\,
            DIN => \N__40058\,
            DOUT => \N__40057\,
            PACKAGEPIN => hsync_wire
        );

    \hsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40059\,
            PADOUT => \N__40058\,
            PADIN => \N__40057\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12935\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40050\,
            DIN => \N__40049\,
            DOUT => \N__40048\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40050\,
            PADOUT => \N__40049\,
            PADIN => \N__40048\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__25805\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40041\,
            DIN => \N__40040\,
            DOUT => \N__40039\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40041\,
            PADOUT => \N__40040\,
            PADIN => \N__40039\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__38012\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40032\,
            DIN => \N__40031\,
            DOUT => \N__40030\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40032\,
            PADOUT => \N__40031\,
            PADIN => \N__40030\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40023\,
            DIN => \N__40022\,
            DOUT => \N__40021\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40023\,
            PADOUT => \N__40022\,
            PADIN => \N__40021\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40014\,
            DIN => \N__40013\,
            DOUT => \N__40012\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40014\,
            PADOUT => \N__40013\,
            PADIN => \N__40012\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__40005\,
            DIN => \N__40004\,
            DOUT => \N__40003\,
            PACKAGEPIN => led_wire(5)
        );

    \led_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__40005\,
            PADOUT => \N__40004\,
            PADIN => \N__40003\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39996\,
            DIN => \N__39995\,
            DOUT => \N__39994\,
            PACKAGEPIN => led_wire(6)
        );

    \led_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39996\,
            PADOUT => \N__39995\,
            PADIN => \N__39994\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__34400\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \led_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39987\,
            DIN => \N__39986\,
            DOUT => \N__39985\,
            PACKAGEPIN => led_wire(7)
        );

    \led_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39987\,
            PADOUT => \N__39986\,
            PADIN => \N__39985\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37913\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_address_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39978\,
            DIN => \N__39977\,
            DOUT => \N__39976\,
            PACKAGEPIN => port_address(0)
        );

    \port_address_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39978\,
            PADOUT => \N__39977\,
            PADIN => \N__39976\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_0,
            DIN1 => OPEN,
            DOUT0 => \N__35858\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15372\
        );

    \port_address_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39969\,
            DIN => \N__39968\,
            DOUT => \N__39967\,
            PACKAGEPIN => port_address(1)
        );

    \port_address_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39969\,
            PADOUT => \N__39968\,
            PADIN => \N__39967\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_1,
            DIN1 => OPEN,
            DOUT0 => \N__35840\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15404\
        );

    \port_address_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39960\,
            DIN => \N__39959\,
            DOUT => \N__39958\,
            PACKAGEPIN => port_address(2)
        );

    \port_address_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39960\,
            PADOUT => \N__39959\,
            PADIN => \N__39958\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_2,
            DIN1 => OPEN,
            DOUT0 => \N__36392\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15362\
        );

    \port_address_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39951\,
            DIN => \N__39950\,
            DOUT => \N__39949\,
            PACKAGEPIN => port_address(3)
        );

    \port_address_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39951\,
            PADOUT => \N__39950\,
            PADIN => \N__39949\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_3,
            DIN1 => OPEN,
            DOUT0 => \N__36368\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15440\
        );

    \port_address_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39942\,
            DIN => \N__39941\,
            DOUT => \N__39940\,
            PACKAGEPIN => port_address(4)
        );

    \port_address_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39942\,
            PADOUT => \N__39941\,
            PADIN => \N__39940\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_4,
            DIN1 => OPEN,
            DOUT0 => \N__36341\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15435\
        );

    \port_address_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39933\,
            DIN => \N__39932\,
            DOUT => \N__39931\,
            PACKAGEPIN => port_address(5)
        );

    \port_address_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39933\,
            PADOUT => \N__39932\,
            PADIN => \N__39931\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_5,
            DIN1 => OPEN,
            DOUT0 => \N__36314\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15424\
        );

    \port_address_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39924\,
            DIN => \N__39923\,
            DOUT => \N__39922\,
            PACKAGEPIN => port_address(6)
        );

    \port_address_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39924\,
            PADOUT => \N__39923\,
            PADIN => \N__39922\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_6,
            DIN1 => OPEN,
            DOUT0 => \N__36287\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15409\
        );

    \port_address_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39915\,
            DIN => \N__39914\,
            DOUT => \N__39913\,
            PACKAGEPIN => port_address(7)
        );

    \port_address_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39915\,
            PADOUT => \N__39914\,
            PADIN => \N__39913\,
            CLOCKENABLE => 'H',
            DIN0 => port_address_in_7,
            DIN1 => OPEN,
            DOUT0 => \N__36257\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15373\
        );

    \port_address_obuft_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39906\,
            DIN => \N__39905\,
            DOUT => \N__39904\,
            PACKAGEPIN => port_address(10)
        );

    \port_address_obuft_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39906\,
            PADOUT => \N__39905\,
            PADIN => \N__39904\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37250\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15364\
        );

    \port_address_obuft_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39897\,
            DIN => \N__39896\,
            DOUT => \N__39895\,
            PACKAGEPIN => port_address(11)
        );

    \port_address_obuft_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39897\,
            PADOUT => \N__39896\,
            PADIN => \N__39895\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37223\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15423\
        );

    \port_address_obuft_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39888\,
            DIN => \N__39887\,
            DOUT => \N__39886\,
            PACKAGEPIN => port_address(12)
        );

    \port_address_obuft_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39888\,
            PADOUT => \N__39887\,
            PADIN => \N__39886\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37190\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15436\
        );

    \port_address_obuft_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39879\,
            DIN => \N__39878\,
            DOUT => \N__39877\,
            PACKAGEPIN => port_address(13)
        );

    \port_address_obuft_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39879\,
            PADOUT => \N__39878\,
            PADIN => \N__39877\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37160\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15425\
        );

    \port_address_obuft_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39870\,
            DIN => \N__39869\,
            DOUT => \N__39868\,
            PACKAGEPIN => port_address(14)
        );

    \port_address_obuft_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39870\,
            PADOUT => \N__39869\,
            PADIN => \N__39868\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37130\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15408\
        );

    \port_address_obuft_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39861\,
            DIN => \N__39860\,
            DOUT => \N__39859\,
            PACKAGEPIN => port_address(15)
        );

    \port_address_obuft_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39861\,
            PADOUT => \N__39860\,
            PADIN => \N__39859\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__37019\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15311\
        );

    \port_address_obuft_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39852\,
            DIN => \N__39851\,
            DOUT => \N__39850\,
            PACKAGEPIN => port_address(8)
        );

    \port_address_obuft_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39852\,
            PADOUT => \N__39851\,
            PADIN => \N__39850\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36227\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15363\
        );

    \port_address_obuft_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39843\,
            DIN => \N__39842\,
            DOUT => \N__39841\,
            PACKAGEPIN => port_address(9)
        );

    \port_address_obuft_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39843\,
            PADOUT => \N__39842\,
            PADIN => \N__39841\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__36197\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15403\
        );

    \port_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39834\,
            DIN => \N__39833\,
            DOUT => \N__39832\,
            PACKAGEPIN => port_clk_wire
        );

    \port_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39834\,
            PADOUT => \N__39833\,
            PADIN => \N__39832\,
            CLOCKENABLE => 'H',
            DIN0 => port_clk_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39825\,
            DIN => \N__39824\,
            DOUT => \N__39823\,
            PACKAGEPIN => port_data_wire(0)
        );

    \port_data_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39825\,
            PADOUT => \N__39824\,
            PADIN => \N__39823\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39816\,
            DIN => \N__39815\,
            DOUT => \N__39814\,
            PACKAGEPIN => port_data_wire(1)
        );

    \port_data_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39816\,
            PADOUT => \N__39815\,
            PADIN => \N__39814\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39807\,
            DIN => \N__39806\,
            DOUT => \N__39805\,
            PACKAGEPIN => port_data_wire(2)
        );

    \port_data_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39807\,
            PADOUT => \N__39806\,
            PADIN => \N__39805\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39798\,
            DIN => \N__39797\,
            DOUT => \N__39796\,
            PACKAGEPIN => port_data_wire(3)
        );

    \port_data_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39798\,
            PADOUT => \N__39797\,
            PADIN => \N__39796\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39789\,
            DIN => \N__39788\,
            DOUT => \N__39787\,
            PACKAGEPIN => port_data_wire(4)
        );

    \port_data_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39789\,
            PADOUT => \N__39788\,
            PADIN => \N__39787\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39780\,
            DIN => \N__39779\,
            DOUT => \N__39778\,
            PACKAGEPIN => port_data_wire(5)
        );

    \port_data_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39780\,
            PADOUT => \N__39779\,
            PADIN => \N__39778\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39771\,
            DIN => \N__39770\,
            DOUT => \N__39769\,
            PACKAGEPIN => port_data_wire(6)
        );

    \port_data_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39771\,
            PADOUT => \N__39770\,
            PADIN => \N__39769\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39762\,
            DIN => \N__39761\,
            DOUT => \N__39760\,
            PACKAGEPIN => port_data_wire(7)
        );

    \port_data_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39762\,
            PADOUT => \N__39761\,
            PADIN => \N__39760\,
            CLOCKENABLE => 'H',
            DIN0 => port_data_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_data_rw_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39753\,
            DIN => \N__39752\,
            DOUT => \N__39751\,
            PACKAGEPIN => port_data_rw_wire
        );

    \port_data_rw_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39753\,
            PADOUT => \N__39752\,
            PADIN => \N__39751\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12716\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_dmab_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39744\,
            DIN => \N__39743\,
            DOUT => \N__39742\,
            PACKAGEPIN => port_dmab_wire
        );

    \port_dmab_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39744\,
            PADOUT => \N__39743\,
            PADIN => \N__39742\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__34177\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_enb_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39735\,
            DIN => \N__39734\,
            DOUT => \N__39733\,
            PACKAGEPIN => port_enb_wire
        );

    \port_enb_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39735\,
            PADOUT => \N__39734\,
            PADIN => \N__39733\,
            CLOCKENABLE => 'H',
            DIN0 => port_enb_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_nmib_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39726\,
            DIN => \N__39725\,
            DOUT => \N__39724\,
            PACKAGEPIN => port_nmib_wire
        );

    \port_nmib_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39726\,
            PADOUT => \N__39725\,
            PADIN => \N__39724\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__26387\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \port_rw_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39717\,
            DIN => \N__39716\,
            DOUT => \N__39715\,
            PACKAGEPIN => port_rw
        );

    \port_rw_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__39717\,
            PADOUT => \N__39716\,
            PADIN => \N__39715\,
            CLOCKENABLE => 'H',
            DIN0 => port_rw_in,
            DIN1 => OPEN,
            DOUT0 => \N__25682\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__15352\
        );

    \rgb_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39708\,
            DIN => \N__39707\,
            DOUT => \N__39706\,
            PACKAGEPIN => rgb_wire(0)
        );

    \rgb_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39708\,
            PADOUT => \N__39707\,
            PADIN => \N__39706\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12890\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39699\,
            DIN => \N__39698\,
            DOUT => \N__39697\,
            PACKAGEPIN => rgb_wire(1)
        );

    \rgb_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39699\,
            PADOUT => \N__39698\,
            PADIN => \N__39697\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12791\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39690\,
            DIN => \N__39689\,
            DOUT => \N__39688\,
            PACKAGEPIN => rgb_wire(2)
        );

    \rgb_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39690\,
            PADOUT => \N__39689\,
            PADIN => \N__39688\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12770\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39681\,
            DIN => \N__39680\,
            DOUT => \N__39679\,
            PACKAGEPIN => rgb_wire(3)
        );

    \rgb_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39681\,
            PADOUT => \N__39680\,
            PADIN => \N__39679\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12809\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39672\,
            DIN => \N__39671\,
            DOUT => \N__39670\,
            PACKAGEPIN => rgb_wire(4)
        );

    \rgb_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39672\,
            PADOUT => \N__39671\,
            PADIN => \N__39670\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12761\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rgb_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39663\,
            DIN => \N__39662\,
            DOUT => \N__39661\,
            PACKAGEPIN => rgb_wire(5)
        );

    \rgb_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39663\,
            PADOUT => \N__39662\,
            PADIN => \N__39661\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12743\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39654\,
            DIN => \N__39653\,
            DOUT => \N__39652\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__39654\,
            PADOUT => \N__39653\,
            PADIN => \N__39652\,
            CLOCKENABLE => 'H',
            DIN0 => rst_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vblank_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39645\,
            DIN => \N__39644\,
            DOUT => \N__39643\,
            PACKAGEPIN => vblank_wire
        );

    \vblank_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39645\,
            PADOUT => \N__39644\,
            PADIN => \N__39643\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__12899\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \vsync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39636\,
            DIN => \N__39635\,
            DOUT => \N__39634\,
            PACKAGEPIN => vsync_wire
        );

    \vsync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__39636\,
            PADOUT => \N__39635\,
            PADIN => \N__39634\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29879\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__9910\ : CascadeMux
    port map (
            O => \N__39617\,
            I => \N__39614\
        );

    \I__9909\ : CascadeBuf
    port map (
            O => \N__39614\,
            I => \N__39611\
        );

    \I__9908\ : CascadeMux
    port map (
            O => \N__39611\,
            I => \N__39608\
        );

    \I__9907\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39604\
        );

    \I__9906\ : InMux
    port map (
            O => \N__39607\,
            I => \N__39601\
        );

    \I__9905\ : LocalMux
    port map (
            O => \N__39604\,
            I => \N__39598\
        );

    \I__9904\ : LocalMux
    port map (
            O => \N__39601\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__39598\,
            I => \M_this_map_address_qZ0Z_6\
        );

    \I__9902\ : InMux
    port map (
            O => \N__39593\,
            I => \un1_M_this_map_address_q_cry_5\
        );

    \I__9901\ : CascadeMux
    port map (
            O => \N__39590\,
            I => \N__39587\
        );

    \I__9900\ : CascadeBuf
    port map (
            O => \N__39587\,
            I => \N__39584\
        );

    \I__9899\ : CascadeMux
    port map (
            O => \N__39584\,
            I => \N__39581\
        );

    \I__9898\ : InMux
    port map (
            O => \N__39581\,
            I => \N__39578\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__39578\,
            I => \N__39574\
        );

    \I__9896\ : InMux
    port map (
            O => \N__39577\,
            I => \N__39571\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__39574\,
            I => \N__39568\
        );

    \I__9894\ : LocalMux
    port map (
            O => \N__39571\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__9893\ : Odrv4
    port map (
            O => \N__39568\,
            I => \M_this_map_address_qZ0Z_7\
        );

    \I__9892\ : InMux
    port map (
            O => \N__39563\,
            I => \un1_M_this_map_address_q_cry_6\
        );

    \I__9891\ : CascadeMux
    port map (
            O => \N__39560\,
            I => \N__39557\
        );

    \I__9890\ : CascadeBuf
    port map (
            O => \N__39557\,
            I => \N__39554\
        );

    \I__9889\ : CascadeMux
    port map (
            O => \N__39554\,
            I => \N__39551\
        );

    \I__9888\ : InMux
    port map (
            O => \N__39551\,
            I => \N__39548\
        );

    \I__9887\ : LocalMux
    port map (
            O => \N__39548\,
            I => \N__39544\
        );

    \I__9886\ : InMux
    port map (
            O => \N__39547\,
            I => \N__39541\
        );

    \I__9885\ : Span4Mux_h
    port map (
            O => \N__39544\,
            I => \N__39538\
        );

    \I__9884\ : LocalMux
    port map (
            O => \N__39541\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__9883\ : Odrv4
    port map (
            O => \N__39538\,
            I => \M_this_map_address_qZ0Z_8\
        );

    \I__9882\ : InMux
    port map (
            O => \N__39533\,
            I => \bfn_26_26_0_\
        );

    \I__9881\ : CascadeMux
    port map (
            O => \N__39530\,
            I => \N__39527\
        );

    \I__9880\ : InMux
    port map (
            O => \N__39527\,
            I => \N__39514\
        );

    \I__9879\ : InMux
    port map (
            O => \N__39526\,
            I => \N__39509\
        );

    \I__9878\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39509\
        );

    \I__9877\ : InMux
    port map (
            O => \N__39524\,
            I => \N__39500\
        );

    \I__9876\ : InMux
    port map (
            O => \N__39523\,
            I => \N__39500\
        );

    \I__9875\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39500\
        );

    \I__9874\ : InMux
    port map (
            O => \N__39521\,
            I => \N__39500\
        );

    \I__9873\ : InMux
    port map (
            O => \N__39520\,
            I => \N__39491\
        );

    \I__9872\ : InMux
    port map (
            O => \N__39519\,
            I => \N__39491\
        );

    \I__9871\ : InMux
    port map (
            O => \N__39518\,
            I => \N__39491\
        );

    \I__9870\ : InMux
    port map (
            O => \N__39517\,
            I => \N__39491\
        );

    \I__9869\ : LocalMux
    port map (
            O => \N__39514\,
            I => \N__39488\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__39509\,
            I => \N__39481\
        );

    \I__9867\ : LocalMux
    port map (
            O => \N__39500\,
            I => \N__39481\
        );

    \I__9866\ : LocalMux
    port map (
            O => \N__39491\,
            I => \N__39481\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__39488\,
            I => \N__39478\
        );

    \I__9864\ : Span4Mux_v
    port map (
            O => \N__39481\,
            I => \N__39475\
        );

    \I__9863\ : Span4Mux_h
    port map (
            O => \N__39478\,
            I => \N__39472\
        );

    \I__9862\ : Span4Mux_h
    port map (
            O => \N__39475\,
            I => \N__39469\
        );

    \I__9861\ : Odrv4
    port map (
            O => \N__39472\,
            I => \N_93\
        );

    \I__9860\ : Odrv4
    port map (
            O => \N__39469\,
            I => \N_93\
        );

    \I__9859\ : InMux
    port map (
            O => \N__39464\,
            I => \un1_M_this_map_address_q_cry_8\
        );

    \I__9858\ : CascadeMux
    port map (
            O => \N__39461\,
            I => \N__39458\
        );

    \I__9857\ : CascadeBuf
    port map (
            O => \N__39458\,
            I => \N__39455\
        );

    \I__9856\ : CascadeMux
    port map (
            O => \N__39455\,
            I => \N__39452\
        );

    \I__9855\ : InMux
    port map (
            O => \N__39452\,
            I => \N__39449\
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39445\
        );

    \I__9853\ : InMux
    port map (
            O => \N__39448\,
            I => \N__39442\
        );

    \I__9852\ : Span4Mux_h
    port map (
            O => \N__39445\,
            I => \N__39439\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__39442\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__9850\ : Odrv4
    port map (
            O => \N__39439\,
            I => \M_this_map_address_qZ0Z_9\
        );

    \I__9849\ : ClkMux
    port map (
            O => \N__39434\,
            I => \N__38969\
        );

    \I__9848\ : ClkMux
    port map (
            O => \N__39433\,
            I => \N__38969\
        );

    \I__9847\ : ClkMux
    port map (
            O => \N__39432\,
            I => \N__38969\
        );

    \I__9846\ : ClkMux
    port map (
            O => \N__39431\,
            I => \N__38969\
        );

    \I__9845\ : ClkMux
    port map (
            O => \N__39430\,
            I => \N__38969\
        );

    \I__9844\ : ClkMux
    port map (
            O => \N__39429\,
            I => \N__38969\
        );

    \I__9843\ : ClkMux
    port map (
            O => \N__39428\,
            I => \N__38969\
        );

    \I__9842\ : ClkMux
    port map (
            O => \N__39427\,
            I => \N__38969\
        );

    \I__9841\ : ClkMux
    port map (
            O => \N__39426\,
            I => \N__38969\
        );

    \I__9840\ : ClkMux
    port map (
            O => \N__39425\,
            I => \N__38969\
        );

    \I__9839\ : ClkMux
    port map (
            O => \N__39424\,
            I => \N__38969\
        );

    \I__9838\ : ClkMux
    port map (
            O => \N__39423\,
            I => \N__38969\
        );

    \I__9837\ : ClkMux
    port map (
            O => \N__39422\,
            I => \N__38969\
        );

    \I__9836\ : ClkMux
    port map (
            O => \N__39421\,
            I => \N__38969\
        );

    \I__9835\ : ClkMux
    port map (
            O => \N__39420\,
            I => \N__38969\
        );

    \I__9834\ : ClkMux
    port map (
            O => \N__39419\,
            I => \N__38969\
        );

    \I__9833\ : ClkMux
    port map (
            O => \N__39418\,
            I => \N__38969\
        );

    \I__9832\ : ClkMux
    port map (
            O => \N__39417\,
            I => \N__38969\
        );

    \I__9831\ : ClkMux
    port map (
            O => \N__39416\,
            I => \N__38969\
        );

    \I__9830\ : ClkMux
    port map (
            O => \N__39415\,
            I => \N__38969\
        );

    \I__9829\ : ClkMux
    port map (
            O => \N__39414\,
            I => \N__38969\
        );

    \I__9828\ : ClkMux
    port map (
            O => \N__39413\,
            I => \N__38969\
        );

    \I__9827\ : ClkMux
    port map (
            O => \N__39412\,
            I => \N__38969\
        );

    \I__9826\ : ClkMux
    port map (
            O => \N__39411\,
            I => \N__38969\
        );

    \I__9825\ : ClkMux
    port map (
            O => \N__39410\,
            I => \N__38969\
        );

    \I__9824\ : ClkMux
    port map (
            O => \N__39409\,
            I => \N__38969\
        );

    \I__9823\ : ClkMux
    port map (
            O => \N__39408\,
            I => \N__38969\
        );

    \I__9822\ : ClkMux
    port map (
            O => \N__39407\,
            I => \N__38969\
        );

    \I__9821\ : ClkMux
    port map (
            O => \N__39406\,
            I => \N__38969\
        );

    \I__9820\ : ClkMux
    port map (
            O => \N__39405\,
            I => \N__38969\
        );

    \I__9819\ : ClkMux
    port map (
            O => \N__39404\,
            I => \N__38969\
        );

    \I__9818\ : ClkMux
    port map (
            O => \N__39403\,
            I => \N__38969\
        );

    \I__9817\ : ClkMux
    port map (
            O => \N__39402\,
            I => \N__38969\
        );

    \I__9816\ : ClkMux
    port map (
            O => \N__39401\,
            I => \N__38969\
        );

    \I__9815\ : ClkMux
    port map (
            O => \N__39400\,
            I => \N__38969\
        );

    \I__9814\ : ClkMux
    port map (
            O => \N__39399\,
            I => \N__38969\
        );

    \I__9813\ : ClkMux
    port map (
            O => \N__39398\,
            I => \N__38969\
        );

    \I__9812\ : ClkMux
    port map (
            O => \N__39397\,
            I => \N__38969\
        );

    \I__9811\ : ClkMux
    port map (
            O => \N__39396\,
            I => \N__38969\
        );

    \I__9810\ : ClkMux
    port map (
            O => \N__39395\,
            I => \N__38969\
        );

    \I__9809\ : ClkMux
    port map (
            O => \N__39394\,
            I => \N__38969\
        );

    \I__9808\ : ClkMux
    port map (
            O => \N__39393\,
            I => \N__38969\
        );

    \I__9807\ : ClkMux
    port map (
            O => \N__39392\,
            I => \N__38969\
        );

    \I__9806\ : ClkMux
    port map (
            O => \N__39391\,
            I => \N__38969\
        );

    \I__9805\ : ClkMux
    port map (
            O => \N__39390\,
            I => \N__38969\
        );

    \I__9804\ : ClkMux
    port map (
            O => \N__39389\,
            I => \N__38969\
        );

    \I__9803\ : ClkMux
    port map (
            O => \N__39388\,
            I => \N__38969\
        );

    \I__9802\ : ClkMux
    port map (
            O => \N__39387\,
            I => \N__38969\
        );

    \I__9801\ : ClkMux
    port map (
            O => \N__39386\,
            I => \N__38969\
        );

    \I__9800\ : ClkMux
    port map (
            O => \N__39385\,
            I => \N__38969\
        );

    \I__9799\ : ClkMux
    port map (
            O => \N__39384\,
            I => \N__38969\
        );

    \I__9798\ : ClkMux
    port map (
            O => \N__39383\,
            I => \N__38969\
        );

    \I__9797\ : ClkMux
    port map (
            O => \N__39382\,
            I => \N__38969\
        );

    \I__9796\ : ClkMux
    port map (
            O => \N__39381\,
            I => \N__38969\
        );

    \I__9795\ : ClkMux
    port map (
            O => \N__39380\,
            I => \N__38969\
        );

    \I__9794\ : ClkMux
    port map (
            O => \N__39379\,
            I => \N__38969\
        );

    \I__9793\ : ClkMux
    port map (
            O => \N__39378\,
            I => \N__38969\
        );

    \I__9792\ : ClkMux
    port map (
            O => \N__39377\,
            I => \N__38969\
        );

    \I__9791\ : ClkMux
    port map (
            O => \N__39376\,
            I => \N__38969\
        );

    \I__9790\ : ClkMux
    port map (
            O => \N__39375\,
            I => \N__38969\
        );

    \I__9789\ : ClkMux
    port map (
            O => \N__39374\,
            I => \N__38969\
        );

    \I__9788\ : ClkMux
    port map (
            O => \N__39373\,
            I => \N__38969\
        );

    \I__9787\ : ClkMux
    port map (
            O => \N__39372\,
            I => \N__38969\
        );

    \I__9786\ : ClkMux
    port map (
            O => \N__39371\,
            I => \N__38969\
        );

    \I__9785\ : ClkMux
    port map (
            O => \N__39370\,
            I => \N__38969\
        );

    \I__9784\ : ClkMux
    port map (
            O => \N__39369\,
            I => \N__38969\
        );

    \I__9783\ : ClkMux
    port map (
            O => \N__39368\,
            I => \N__38969\
        );

    \I__9782\ : ClkMux
    port map (
            O => \N__39367\,
            I => \N__38969\
        );

    \I__9781\ : ClkMux
    port map (
            O => \N__39366\,
            I => \N__38969\
        );

    \I__9780\ : ClkMux
    port map (
            O => \N__39365\,
            I => \N__38969\
        );

    \I__9779\ : ClkMux
    port map (
            O => \N__39364\,
            I => \N__38969\
        );

    \I__9778\ : ClkMux
    port map (
            O => \N__39363\,
            I => \N__38969\
        );

    \I__9777\ : ClkMux
    port map (
            O => \N__39362\,
            I => \N__38969\
        );

    \I__9776\ : ClkMux
    port map (
            O => \N__39361\,
            I => \N__38969\
        );

    \I__9775\ : ClkMux
    port map (
            O => \N__39360\,
            I => \N__38969\
        );

    \I__9774\ : ClkMux
    port map (
            O => \N__39359\,
            I => \N__38969\
        );

    \I__9773\ : ClkMux
    port map (
            O => \N__39358\,
            I => \N__38969\
        );

    \I__9772\ : ClkMux
    port map (
            O => \N__39357\,
            I => \N__38969\
        );

    \I__9771\ : ClkMux
    port map (
            O => \N__39356\,
            I => \N__38969\
        );

    \I__9770\ : ClkMux
    port map (
            O => \N__39355\,
            I => \N__38969\
        );

    \I__9769\ : ClkMux
    port map (
            O => \N__39354\,
            I => \N__38969\
        );

    \I__9768\ : ClkMux
    port map (
            O => \N__39353\,
            I => \N__38969\
        );

    \I__9767\ : ClkMux
    port map (
            O => \N__39352\,
            I => \N__38969\
        );

    \I__9766\ : ClkMux
    port map (
            O => \N__39351\,
            I => \N__38969\
        );

    \I__9765\ : ClkMux
    port map (
            O => \N__39350\,
            I => \N__38969\
        );

    \I__9764\ : ClkMux
    port map (
            O => \N__39349\,
            I => \N__38969\
        );

    \I__9763\ : ClkMux
    port map (
            O => \N__39348\,
            I => \N__38969\
        );

    \I__9762\ : ClkMux
    port map (
            O => \N__39347\,
            I => \N__38969\
        );

    \I__9761\ : ClkMux
    port map (
            O => \N__39346\,
            I => \N__38969\
        );

    \I__9760\ : ClkMux
    port map (
            O => \N__39345\,
            I => \N__38969\
        );

    \I__9759\ : ClkMux
    port map (
            O => \N__39344\,
            I => \N__38969\
        );

    \I__9758\ : ClkMux
    port map (
            O => \N__39343\,
            I => \N__38969\
        );

    \I__9757\ : ClkMux
    port map (
            O => \N__39342\,
            I => \N__38969\
        );

    \I__9756\ : ClkMux
    port map (
            O => \N__39341\,
            I => \N__38969\
        );

    \I__9755\ : ClkMux
    port map (
            O => \N__39340\,
            I => \N__38969\
        );

    \I__9754\ : ClkMux
    port map (
            O => \N__39339\,
            I => \N__38969\
        );

    \I__9753\ : ClkMux
    port map (
            O => \N__39338\,
            I => \N__38969\
        );

    \I__9752\ : ClkMux
    port map (
            O => \N__39337\,
            I => \N__38969\
        );

    \I__9751\ : ClkMux
    port map (
            O => \N__39336\,
            I => \N__38969\
        );

    \I__9750\ : ClkMux
    port map (
            O => \N__39335\,
            I => \N__38969\
        );

    \I__9749\ : ClkMux
    port map (
            O => \N__39334\,
            I => \N__38969\
        );

    \I__9748\ : ClkMux
    port map (
            O => \N__39333\,
            I => \N__38969\
        );

    \I__9747\ : ClkMux
    port map (
            O => \N__39332\,
            I => \N__38969\
        );

    \I__9746\ : ClkMux
    port map (
            O => \N__39331\,
            I => \N__38969\
        );

    \I__9745\ : ClkMux
    port map (
            O => \N__39330\,
            I => \N__38969\
        );

    \I__9744\ : ClkMux
    port map (
            O => \N__39329\,
            I => \N__38969\
        );

    \I__9743\ : ClkMux
    port map (
            O => \N__39328\,
            I => \N__38969\
        );

    \I__9742\ : ClkMux
    port map (
            O => \N__39327\,
            I => \N__38969\
        );

    \I__9741\ : ClkMux
    port map (
            O => \N__39326\,
            I => \N__38969\
        );

    \I__9740\ : ClkMux
    port map (
            O => \N__39325\,
            I => \N__38969\
        );

    \I__9739\ : ClkMux
    port map (
            O => \N__39324\,
            I => \N__38969\
        );

    \I__9738\ : ClkMux
    port map (
            O => \N__39323\,
            I => \N__38969\
        );

    \I__9737\ : ClkMux
    port map (
            O => \N__39322\,
            I => \N__38969\
        );

    \I__9736\ : ClkMux
    port map (
            O => \N__39321\,
            I => \N__38969\
        );

    \I__9735\ : ClkMux
    port map (
            O => \N__39320\,
            I => \N__38969\
        );

    \I__9734\ : ClkMux
    port map (
            O => \N__39319\,
            I => \N__38969\
        );

    \I__9733\ : ClkMux
    port map (
            O => \N__39318\,
            I => \N__38969\
        );

    \I__9732\ : ClkMux
    port map (
            O => \N__39317\,
            I => \N__38969\
        );

    \I__9731\ : ClkMux
    port map (
            O => \N__39316\,
            I => \N__38969\
        );

    \I__9730\ : ClkMux
    port map (
            O => \N__39315\,
            I => \N__38969\
        );

    \I__9729\ : ClkMux
    port map (
            O => \N__39314\,
            I => \N__38969\
        );

    \I__9728\ : ClkMux
    port map (
            O => \N__39313\,
            I => \N__38969\
        );

    \I__9727\ : ClkMux
    port map (
            O => \N__39312\,
            I => \N__38969\
        );

    \I__9726\ : ClkMux
    port map (
            O => \N__39311\,
            I => \N__38969\
        );

    \I__9725\ : ClkMux
    port map (
            O => \N__39310\,
            I => \N__38969\
        );

    \I__9724\ : ClkMux
    port map (
            O => \N__39309\,
            I => \N__38969\
        );

    \I__9723\ : ClkMux
    port map (
            O => \N__39308\,
            I => \N__38969\
        );

    \I__9722\ : ClkMux
    port map (
            O => \N__39307\,
            I => \N__38969\
        );

    \I__9721\ : ClkMux
    port map (
            O => \N__39306\,
            I => \N__38969\
        );

    \I__9720\ : ClkMux
    port map (
            O => \N__39305\,
            I => \N__38969\
        );

    \I__9719\ : ClkMux
    port map (
            O => \N__39304\,
            I => \N__38969\
        );

    \I__9718\ : ClkMux
    port map (
            O => \N__39303\,
            I => \N__38969\
        );

    \I__9717\ : ClkMux
    port map (
            O => \N__39302\,
            I => \N__38969\
        );

    \I__9716\ : ClkMux
    port map (
            O => \N__39301\,
            I => \N__38969\
        );

    \I__9715\ : ClkMux
    port map (
            O => \N__39300\,
            I => \N__38969\
        );

    \I__9714\ : ClkMux
    port map (
            O => \N__39299\,
            I => \N__38969\
        );

    \I__9713\ : ClkMux
    port map (
            O => \N__39298\,
            I => \N__38969\
        );

    \I__9712\ : ClkMux
    port map (
            O => \N__39297\,
            I => \N__38969\
        );

    \I__9711\ : ClkMux
    port map (
            O => \N__39296\,
            I => \N__38969\
        );

    \I__9710\ : ClkMux
    port map (
            O => \N__39295\,
            I => \N__38969\
        );

    \I__9709\ : ClkMux
    port map (
            O => \N__39294\,
            I => \N__38969\
        );

    \I__9708\ : ClkMux
    port map (
            O => \N__39293\,
            I => \N__38969\
        );

    \I__9707\ : ClkMux
    port map (
            O => \N__39292\,
            I => \N__38969\
        );

    \I__9706\ : ClkMux
    port map (
            O => \N__39291\,
            I => \N__38969\
        );

    \I__9705\ : ClkMux
    port map (
            O => \N__39290\,
            I => \N__38969\
        );

    \I__9704\ : ClkMux
    port map (
            O => \N__39289\,
            I => \N__38969\
        );

    \I__9703\ : ClkMux
    port map (
            O => \N__39288\,
            I => \N__38969\
        );

    \I__9702\ : ClkMux
    port map (
            O => \N__39287\,
            I => \N__38969\
        );

    \I__9701\ : ClkMux
    port map (
            O => \N__39286\,
            I => \N__38969\
        );

    \I__9700\ : ClkMux
    port map (
            O => \N__39285\,
            I => \N__38969\
        );

    \I__9699\ : ClkMux
    port map (
            O => \N__39284\,
            I => \N__38969\
        );

    \I__9698\ : ClkMux
    port map (
            O => \N__39283\,
            I => \N__38969\
        );

    \I__9697\ : ClkMux
    port map (
            O => \N__39282\,
            I => \N__38969\
        );

    \I__9696\ : ClkMux
    port map (
            O => \N__39281\,
            I => \N__38969\
        );

    \I__9695\ : ClkMux
    port map (
            O => \N__39280\,
            I => \N__38969\
        );

    \I__9694\ : GlobalMux
    port map (
            O => \N__38969\,
            I => \N__38966\
        );

    \I__9693\ : gio2CtrlBuf
    port map (
            O => \N__38966\,
            I => clk_0_c_g
        );

    \I__9692\ : SRMux
    port map (
            O => \N__38963\,
            I => \N__38924\
        );

    \I__9691\ : SRMux
    port map (
            O => \N__38962\,
            I => \N__38924\
        );

    \I__9690\ : SRMux
    port map (
            O => \N__38961\,
            I => \N__38924\
        );

    \I__9689\ : SRMux
    port map (
            O => \N__38960\,
            I => \N__38924\
        );

    \I__9688\ : SRMux
    port map (
            O => \N__38959\,
            I => \N__38924\
        );

    \I__9687\ : SRMux
    port map (
            O => \N__38958\,
            I => \N__38924\
        );

    \I__9686\ : SRMux
    port map (
            O => \N__38957\,
            I => \N__38924\
        );

    \I__9685\ : SRMux
    port map (
            O => \N__38956\,
            I => \N__38924\
        );

    \I__9684\ : SRMux
    port map (
            O => \N__38955\,
            I => \N__38924\
        );

    \I__9683\ : SRMux
    port map (
            O => \N__38954\,
            I => \N__38924\
        );

    \I__9682\ : SRMux
    port map (
            O => \N__38953\,
            I => \N__38924\
        );

    \I__9681\ : SRMux
    port map (
            O => \N__38952\,
            I => \N__38924\
        );

    \I__9680\ : SRMux
    port map (
            O => \N__38951\,
            I => \N__38924\
        );

    \I__9679\ : GlobalMux
    port map (
            O => \N__38924\,
            I => \N__38921\
        );

    \I__9678\ : gio2CtrlBuf
    port map (
            O => \N__38921\,
            I => \N_527_g\
        );

    \I__9677\ : InMux
    port map (
            O => \N__38918\,
            I => \N__38914\
        );

    \I__9676\ : InMux
    port map (
            O => \N__38917\,
            I => \N__38911\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__38914\,
            I => \N__38904\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__38911\,
            I => \N__38904\
        );

    \I__9673\ : InMux
    port map (
            O => \N__38910\,
            I => \N__38900\
        );

    \I__9672\ : CascadeMux
    port map (
            O => \N__38909\,
            I => \N__38897\
        );

    \I__9671\ : Span4Mux_v
    port map (
            O => \N__38904\,
            I => \N__38891\
        );

    \I__9670\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38887\
        );

    \I__9669\ : LocalMux
    port map (
            O => \N__38900\,
            I => \N__38883\
        );

    \I__9668\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38880\
        );

    \I__9667\ : CascadeMux
    port map (
            O => \N__38896\,
            I => \N__38877\
        );

    \I__9666\ : InMux
    port map (
            O => \N__38895\,
            I => \N__38874\
        );

    \I__9665\ : InMux
    port map (
            O => \N__38894\,
            I => \N__38871\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__38891\,
            I => \N__38868\
        );

    \I__9663\ : InMux
    port map (
            O => \N__38890\,
            I => \N__38865\
        );

    \I__9662\ : LocalMux
    port map (
            O => \N__38887\,
            I => \N__38862\
        );

    \I__9661\ : InMux
    port map (
            O => \N__38886\,
            I => \N__38859\
        );

    \I__9660\ : Span4Mux_v
    port map (
            O => \N__38883\,
            I => \N__38856\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__38880\,
            I => \N__38853\
        );

    \I__9658\ : InMux
    port map (
            O => \N__38877\,
            I => \N__38850\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__38874\,
            I => \N__38845\
        );

    \I__9656\ : LocalMux
    port map (
            O => \N__38871\,
            I => \N__38845\
        );

    \I__9655\ : Span4Mux_v
    port map (
            O => \N__38868\,
            I => \N__38842\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__38865\,
            I => \N__38839\
        );

    \I__9653\ : Span4Mux_v
    port map (
            O => \N__38862\,
            I => \N__38836\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__38859\,
            I => \N__38833\
        );

    \I__9651\ : Span4Mux_h
    port map (
            O => \N__38856\,
            I => \N__38828\
        );

    \I__9650\ : Span4Mux_v
    port map (
            O => \N__38853\,
            I => \N__38828\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__38850\,
            I => \N__38825\
        );

    \I__9648\ : Span12Mux_h
    port map (
            O => \N__38845\,
            I => \N__38822\
        );

    \I__9647\ : Span4Mux_v
    port map (
            O => \N__38842\,
            I => \N__38817\
        );

    \I__9646\ : Span4Mux_v
    port map (
            O => \N__38839\,
            I => \N__38817\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__38836\,
            I => \N__38812\
        );

    \I__9644\ : Span4Mux_v
    port map (
            O => \N__38833\,
            I => \N__38812\
        );

    \I__9643\ : Span4Mux_h
    port map (
            O => \N__38828\,
            I => \N__38807\
        );

    \I__9642\ : Span4Mux_v
    port map (
            O => \N__38825\,
            I => \N__38807\
        );

    \I__9641\ : Span12Mux_h
    port map (
            O => \N__38822\,
            I => \N__38804\
        );

    \I__9640\ : Sp12to4
    port map (
            O => \N__38817\,
            I => \N__38801\
        );

    \I__9639\ : Span4Mux_v
    port map (
            O => \N__38812\,
            I => \N__38796\
        );

    \I__9638\ : Span4Mux_h
    port map (
            O => \N__38807\,
            I => \N__38796\
        );

    \I__9637\ : Span12Mux_v
    port map (
            O => \N__38804\,
            I => \N__38793\
        );

    \I__9636\ : Span12Mux_h
    port map (
            O => \N__38801\,
            I => \N__38790\
        );

    \I__9635\ : Span4Mux_h
    port map (
            O => \N__38796\,
            I => \N__38787\
        );

    \I__9634\ : Odrv12
    port map (
            O => \N__38793\,
            I => port_data_c_5
        );

    \I__9633\ : Odrv12
    port map (
            O => \N__38790\,
            I => port_data_c_5
        );

    \I__9632\ : Odrv4
    port map (
            O => \N__38787\,
            I => port_data_c_5
        );

    \I__9631\ : InMux
    port map (
            O => \N__38780\,
            I => \N__38777\
        );

    \I__9630\ : LocalMux
    port map (
            O => \N__38777\,
            I => \M_this_map_ram_write_data_5\
        );

    \I__9629\ : InMux
    port map (
            O => \N__38774\,
            I => \N__38770\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__38773\,
            I => \N__38765\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__38770\,
            I => \N__38762\
        );

    \I__9626\ : InMux
    port map (
            O => \N__38769\,
            I => \N__38756\
        );

    \I__9625\ : InMux
    port map (
            O => \N__38768\,
            I => \N__38753\
        );

    \I__9624\ : InMux
    port map (
            O => \N__38765\,
            I => \N__38750\
        );

    \I__9623\ : Span4Mux_v
    port map (
            O => \N__38762\,
            I => \N__38747\
        );

    \I__9622\ : InMux
    port map (
            O => \N__38761\,
            I => \N__38744\
        );

    \I__9621\ : InMux
    port map (
            O => \N__38760\,
            I => \N__38741\
        );

    \I__9620\ : InMux
    port map (
            O => \N__38759\,
            I => \N__38738\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__38756\,
            I => \N__38734\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__38753\,
            I => \N__38731\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__38750\,
            I => \N__38726\
        );

    \I__9616\ : Span4Mux_v
    port map (
            O => \N__38747\,
            I => \N__38723\
        );

    \I__9615\ : LocalMux
    port map (
            O => \N__38744\,
            I => \N__38720\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__38741\,
            I => \N__38715\
        );

    \I__9613\ : LocalMux
    port map (
            O => \N__38738\,
            I => \N__38715\
        );

    \I__9612\ : CascadeMux
    port map (
            O => \N__38737\,
            I => \N__38712\
        );

    \I__9611\ : Span4Mux_h
    port map (
            O => \N__38734\,
            I => \N__38709\
        );

    \I__9610\ : Span4Mux_h
    port map (
            O => \N__38731\,
            I => \N__38706\
        );

    \I__9609\ : InMux
    port map (
            O => \N__38730\,
            I => \N__38703\
        );

    \I__9608\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38700\
        );

    \I__9607\ : Span4Mux_v
    port map (
            O => \N__38726\,
            I => \N__38697\
        );

    \I__9606\ : Span4Mux_v
    port map (
            O => \N__38723\,
            I => \N__38694\
        );

    \I__9605\ : Span4Mux_v
    port map (
            O => \N__38720\,
            I => \N__38689\
        );

    \I__9604\ : Span4Mux_h
    port map (
            O => \N__38715\,
            I => \N__38689\
        );

    \I__9603\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38686\
        );

    \I__9602\ : Sp12to4
    port map (
            O => \N__38709\,
            I => \N__38681\
        );

    \I__9601\ : Sp12to4
    port map (
            O => \N__38706\,
            I => \N__38681\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38676\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38676\
        );

    \I__9598\ : Span4Mux_v
    port map (
            O => \N__38697\,
            I => \N__38667\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__38694\,
            I => \N__38667\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__38689\,
            I => \N__38667\
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__38686\,
            I => \N__38667\
        );

    \I__9594\ : Span12Mux_s10_v
    port map (
            O => \N__38681\,
            I => \N__38664\
        );

    \I__9593\ : Span12Mux_s10_v
    port map (
            O => \N__38676\,
            I => \N__38661\
        );

    \I__9592\ : Span4Mux_v
    port map (
            O => \N__38667\,
            I => \N__38658\
        );

    \I__9591\ : Span12Mux_v
    port map (
            O => \N__38664\,
            I => \N__38655\
        );

    \I__9590\ : Span12Mux_v
    port map (
            O => \N__38661\,
            I => \N__38652\
        );

    \I__9589\ : Span4Mux_v
    port map (
            O => \N__38658\,
            I => \N__38649\
        );

    \I__9588\ : Span12Mux_h
    port map (
            O => \N__38655\,
            I => \N__38646\
        );

    \I__9587\ : Span12Mux_h
    port map (
            O => \N__38652\,
            I => \N__38641\
        );

    \I__9586\ : Sp12to4
    port map (
            O => \N__38649\,
            I => \N__38641\
        );

    \I__9585\ : Odrv12
    port map (
            O => \N__38646\,
            I => port_data_c_7
        );

    \I__9584\ : Odrv12
    port map (
            O => \N__38641\,
            I => port_data_c_7
        );

    \I__9583\ : InMux
    port map (
            O => \N__38636\,
            I => \N__38633\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__38633\,
            I => \M_this_map_ram_write_data_7\
        );

    \I__9581\ : CEMux
    port map (
            O => \N__38630\,
            I => \N__38621\
        );

    \I__9580\ : InMux
    port map (
            O => \N__38629\,
            I => \N__38609\
        );

    \I__9579\ : InMux
    port map (
            O => \N__38628\,
            I => \N__38609\
        );

    \I__9578\ : InMux
    port map (
            O => \N__38627\,
            I => \N__38609\
        );

    \I__9577\ : InMux
    port map (
            O => \N__38626\,
            I => \N__38609\
        );

    \I__9576\ : CEMux
    port map (
            O => \N__38625\,
            I => \N__38606\
        );

    \I__9575\ : InMux
    port map (
            O => \N__38624\,
            I => \N__38603\
        );

    \I__9574\ : LocalMux
    port map (
            O => \N__38621\,
            I => \N__38599\
        );

    \I__9573\ : InMux
    port map (
            O => \N__38620\,
            I => \N__38596\
        );

    \I__9572\ : InMux
    port map (
            O => \N__38619\,
            I => \N__38591\
        );

    \I__9571\ : InMux
    port map (
            O => \N__38618\,
            I => \N__38591\
        );

    \I__9570\ : LocalMux
    port map (
            O => \N__38609\,
            I => \N__38588\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__38606\,
            I => \N__38584\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__38603\,
            I => \N__38581\
        );

    \I__9567\ : CascadeMux
    port map (
            O => \N__38602\,
            I => \N__38578\
        );

    \I__9566\ : Span4Mux_h
    port map (
            O => \N__38599\,
            I => \N__38573\
        );

    \I__9565\ : LocalMux
    port map (
            O => \N__38596\,
            I => \N__38573\
        );

    \I__9564\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38570\
        );

    \I__9563\ : Span4Mux_h
    port map (
            O => \N__38588\,
            I => \N__38567\
        );

    \I__9562\ : InMux
    port map (
            O => \N__38587\,
            I => \N__38564\
        );

    \I__9561\ : Span4Mux_v
    port map (
            O => \N__38584\,
            I => \N__38559\
        );

    \I__9560\ : Span4Mux_h
    port map (
            O => \N__38581\,
            I => \N__38559\
        );

    \I__9559\ : InMux
    port map (
            O => \N__38578\,
            I => \N__38556\
        );

    \I__9558\ : Span4Mux_v
    port map (
            O => \N__38573\,
            I => \N__38553\
        );

    \I__9557\ : Span4Mux_v
    port map (
            O => \N__38570\,
            I => \N__38550\
        );

    \I__9556\ : Span4Mux_v
    port map (
            O => \N__38567\,
            I => \N__38547\
        );

    \I__9555\ : LocalMux
    port map (
            O => \N__38564\,
            I => \N__38540\
        );

    \I__9554\ : Sp12to4
    port map (
            O => \N__38559\,
            I => \N__38540\
        );

    \I__9553\ : LocalMux
    port map (
            O => \N__38556\,
            I => \N__38540\
        );

    \I__9552\ : Span4Mux_h
    port map (
            O => \N__38553\,
            I => \N__38537\
        );

    \I__9551\ : Sp12to4
    port map (
            O => \N__38550\,
            I => \N__38530\
        );

    \I__9550\ : Sp12to4
    port map (
            O => \N__38547\,
            I => \N__38530\
        );

    \I__9549\ : Span12Mux_v
    port map (
            O => \N__38540\,
            I => \N__38530\
        );

    \I__9548\ : Span4Mux_h
    port map (
            O => \N__38537\,
            I => \N__38527\
        );

    \I__9547\ : Span12Mux_h
    port map (
            O => \N__38530\,
            I => \N__38524\
        );

    \I__9546\ : Odrv4
    port map (
            O => \N__38527\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__9545\ : Odrv12
    port map (
            O => \N__38524\,
            I => \M_this_state_d_0_sqmuxa\
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__38519\,
            I => \N__38516\
        );

    \I__9543\ : CascadeBuf
    port map (
            O => \N__38516\,
            I => \N__38513\
        );

    \I__9542\ : CascadeMux
    port map (
            O => \N__38513\,
            I => \N__38510\
        );

    \I__9541\ : InMux
    port map (
            O => \N__38510\,
            I => \N__38506\
        );

    \I__9540\ : InMux
    port map (
            O => \N__38509\,
            I => \N__38503\
        );

    \I__9539\ : LocalMux
    port map (
            O => \N__38506\,
            I => \N__38500\
        );

    \I__9538\ : LocalMux
    port map (
            O => \N__38503\,
            I => \N__38495\
        );

    \I__9537\ : Span4Mux_v
    port map (
            O => \N__38500\,
            I => \N__38495\
        );

    \I__9536\ : Odrv4
    port map (
            O => \N__38495\,
            I => \M_this_map_address_qZ0Z_0\
        );

    \I__9535\ : CascadeMux
    port map (
            O => \N__38492\,
            I => \N__38489\
        );

    \I__9534\ : CascadeBuf
    port map (
            O => \N__38489\,
            I => \N__38486\
        );

    \I__9533\ : CascadeMux
    port map (
            O => \N__38486\,
            I => \N__38483\
        );

    \I__9532\ : InMux
    port map (
            O => \N__38483\,
            I => \N__38480\
        );

    \I__9531\ : LocalMux
    port map (
            O => \N__38480\,
            I => \N__38476\
        );

    \I__9530\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38473\
        );

    \I__9529\ : Span4Mux_v
    port map (
            O => \N__38476\,
            I => \N__38470\
        );

    \I__9528\ : LocalMux
    port map (
            O => \N__38473\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9527\ : Odrv4
    port map (
            O => \N__38470\,
            I => \M_this_map_address_qZ0Z_1\
        );

    \I__9526\ : InMux
    port map (
            O => \N__38465\,
            I => \un1_M_this_map_address_q_cry_0\
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__38462\,
            I => \N__38459\
        );

    \I__9524\ : CascadeBuf
    port map (
            O => \N__38459\,
            I => \N__38456\
        );

    \I__9523\ : CascadeMux
    port map (
            O => \N__38456\,
            I => \N__38453\
        );

    \I__9522\ : InMux
    port map (
            O => \N__38453\,
            I => \N__38450\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38446\
        );

    \I__9520\ : InMux
    port map (
            O => \N__38449\,
            I => \N__38443\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__38446\,
            I => \N__38440\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__38443\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__9517\ : Odrv4
    port map (
            O => \N__38440\,
            I => \M_this_map_address_qZ0Z_2\
        );

    \I__9516\ : InMux
    port map (
            O => \N__38435\,
            I => \un1_M_this_map_address_q_cry_1\
        );

    \I__9515\ : CascadeMux
    port map (
            O => \N__38432\,
            I => \N__38429\
        );

    \I__9514\ : CascadeBuf
    port map (
            O => \N__38429\,
            I => \N__38426\
        );

    \I__9513\ : CascadeMux
    port map (
            O => \N__38426\,
            I => \N__38423\
        );

    \I__9512\ : InMux
    port map (
            O => \N__38423\,
            I => \N__38419\
        );

    \I__9511\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38416\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__38419\,
            I => \N__38413\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__38416\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__9508\ : Odrv4
    port map (
            O => \N__38413\,
            I => \M_this_map_address_qZ0Z_3\
        );

    \I__9507\ : InMux
    port map (
            O => \N__38408\,
            I => \un1_M_this_map_address_q_cry_2\
        );

    \I__9506\ : CascadeMux
    port map (
            O => \N__38405\,
            I => \N__38402\
        );

    \I__9505\ : CascadeBuf
    port map (
            O => \N__38402\,
            I => \N__38399\
        );

    \I__9504\ : CascadeMux
    port map (
            O => \N__38399\,
            I => \N__38396\
        );

    \I__9503\ : InMux
    port map (
            O => \N__38396\,
            I => \N__38393\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38389\
        );

    \I__9501\ : InMux
    port map (
            O => \N__38392\,
            I => \N__38386\
        );

    \I__9500\ : Span4Mux_h
    port map (
            O => \N__38389\,
            I => \N__38383\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__38386\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__9498\ : Odrv4
    port map (
            O => \N__38383\,
            I => \M_this_map_address_qZ0Z_4\
        );

    \I__9497\ : InMux
    port map (
            O => \N__38378\,
            I => \un1_M_this_map_address_q_cry_3\
        );

    \I__9496\ : CascadeMux
    port map (
            O => \N__38375\,
            I => \N__38372\
        );

    \I__9495\ : CascadeBuf
    port map (
            O => \N__38372\,
            I => \N__38369\
        );

    \I__9494\ : CascadeMux
    port map (
            O => \N__38369\,
            I => \N__38366\
        );

    \I__9493\ : InMux
    port map (
            O => \N__38366\,
            I => \N__38362\
        );

    \I__9492\ : InMux
    port map (
            O => \N__38365\,
            I => \N__38359\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__38362\,
            I => \N__38356\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__38359\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__38356\,
            I => \M_this_map_address_qZ0Z_5\
        );

    \I__9488\ : InMux
    port map (
            O => \N__38351\,
            I => \un1_M_this_map_address_q_cry_4\
        );

    \I__9487\ : InMux
    port map (
            O => \N__38348\,
            I => \N__38340\
        );

    \I__9486\ : InMux
    port map (
            O => \N__38347\,
            I => \N__38335\
        );

    \I__9485\ : InMux
    port map (
            O => \N__38346\,
            I => \N__38335\
        );

    \I__9484\ : InMux
    port map (
            O => \N__38345\,
            I => \N__38329\
        );

    \I__9483\ : InMux
    port map (
            O => \N__38344\,
            I => \N__38329\
        );

    \I__9482\ : InMux
    port map (
            O => \N__38343\,
            I => \N__38326\
        );

    \I__9481\ : LocalMux
    port map (
            O => \N__38340\,
            I => \N__38323\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__38335\,
            I => \N__38320\
        );

    \I__9479\ : InMux
    port map (
            O => \N__38334\,
            I => \N__38317\
        );

    \I__9478\ : LocalMux
    port map (
            O => \N__38329\,
            I => \N__38312\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__38326\,
            I => \N__38312\
        );

    \I__9476\ : Span4Mux_h
    port map (
            O => \N__38323\,
            I => \N__38309\
        );

    \I__9475\ : Span4Mux_v
    port map (
            O => \N__38320\,
            I => \N__38301\
        );

    \I__9474\ : LocalMux
    port map (
            O => \N__38317\,
            I => \N__38301\
        );

    \I__9473\ : Span4Mux_v
    port map (
            O => \N__38312\,
            I => \N__38301\
        );

    \I__9472\ : Span4Mux_v
    port map (
            O => \N__38309\,
            I => \N__38298\
        );

    \I__9471\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38295\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__38301\,
            I => \N__38292\
        );

    \I__9469\ : Odrv4
    port map (
            O => \N__38298\,
            I => \N_930\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__38295\,
            I => \N_930\
        );

    \I__9467\ : Odrv4
    port map (
            O => \N__38292\,
            I => \N_930\
        );

    \I__9466\ : InMux
    port map (
            O => \N__38285\,
            I => \N__38274\
        );

    \I__9465\ : InMux
    port map (
            O => \N__38284\,
            I => \N__38271\
        );

    \I__9464\ : InMux
    port map (
            O => \N__38283\,
            I => \N__38268\
        );

    \I__9463\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38264\
        );

    \I__9462\ : InMux
    port map (
            O => \N__38281\,
            I => \N__38261\
        );

    \I__9461\ : InMux
    port map (
            O => \N__38280\,
            I => \N__38258\
        );

    \I__9460\ : InMux
    port map (
            O => \N__38279\,
            I => \N__38255\
        );

    \I__9459\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38252\
        );

    \I__9458\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38249\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__38274\,
            I => \N__38244\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__38271\,
            I => \N__38244\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38241\
        );

    \I__9454\ : InMux
    port map (
            O => \N__38267\,
            I => \N__38238\
        );

    \I__9453\ : LocalMux
    port map (
            O => \N__38264\,
            I => \N__38235\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__38261\,
            I => \N__38230\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__38258\,
            I => \N__38230\
        );

    \I__9450\ : LocalMux
    port map (
            O => \N__38255\,
            I => \N__38222\
        );

    \I__9449\ : LocalMux
    port map (
            O => \N__38252\,
            I => \N__38222\
        );

    \I__9448\ : LocalMux
    port map (
            O => \N__38249\,
            I => \N__38219\
        );

    \I__9447\ : Span4Mux_v
    port map (
            O => \N__38244\,
            I => \N__38214\
        );

    \I__9446\ : Span4Mux_v
    port map (
            O => \N__38241\,
            I => \N__38214\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__38238\,
            I => \N__38211\
        );

    \I__9444\ : Span4Mux_v
    port map (
            O => \N__38235\,
            I => \N__38206\
        );

    \I__9443\ : Span4Mux_h
    port map (
            O => \N__38230\,
            I => \N__38206\
        );

    \I__9442\ : InMux
    port map (
            O => \N__38229\,
            I => \N__38203\
        );

    \I__9441\ : InMux
    port map (
            O => \N__38228\,
            I => \N__38198\
        );

    \I__9440\ : InMux
    port map (
            O => \N__38227\,
            I => \N__38198\
        );

    \I__9439\ : Span12Mux_h
    port map (
            O => \N__38222\,
            I => \N__38195\
        );

    \I__9438\ : Span4Mux_v
    port map (
            O => \N__38219\,
            I => \N__38192\
        );

    \I__9437\ : Span4Mux_h
    port map (
            O => \N__38214\,
            I => \N__38185\
        );

    \I__9436\ : Span4Mux_v
    port map (
            O => \N__38211\,
            I => \N__38185\
        );

    \I__9435\ : Span4Mux_v
    port map (
            O => \N__38206\,
            I => \N__38185\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__38203\,
            I => \N__38180\
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__38198\,
            I => \N__38180\
        );

    \I__9432\ : Odrv12
    port map (
            O => \N__38195\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__9431\ : Odrv4
    port map (
            O => \N__38192\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__9430\ : Odrv4
    port map (
            O => \N__38185\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__9429\ : Odrv12
    port map (
            O => \N__38180\,
            I => \M_this_state_qZ0Z_9\
        );

    \I__9428\ : InMux
    port map (
            O => \N__38171\,
            I => \N__38168\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__38168\,
            I => \N__38165\
        );

    \I__9426\ : Span4Mux_h
    port map (
            O => \N__38165\,
            I => \N__38161\
        );

    \I__9425\ : InMux
    port map (
            O => \N__38164\,
            I => \N__38156\
        );

    \I__9424\ : Span4Mux_h
    port map (
            O => \N__38161\,
            I => \N__38153\
        );

    \I__9423\ : InMux
    port map (
            O => \N__38160\,
            I => \N__38148\
        );

    \I__9422\ : InMux
    port map (
            O => \N__38159\,
            I => \N__38148\
        );

    \I__9421\ : LocalMux
    port map (
            O => \N__38156\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9420\ : Odrv4
    port map (
            O => \N__38153\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9419\ : LocalMux
    port map (
            O => \N__38148\,
            I => \M_this_state_qZ0Z_4\
        );

    \I__9418\ : CascadeMux
    port map (
            O => \N__38141\,
            I => \N__38138\
        );

    \I__9417\ : InMux
    port map (
            O => \N__38138\,
            I => \N__38135\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__38135\,
            I => \N__38132\
        );

    \I__9415\ : Odrv4
    port map (
            O => \N__38132\,
            I => \this_start_data_delay.N_332\
        );

    \I__9414\ : InMux
    port map (
            O => \N__38129\,
            I => \N__38124\
        );

    \I__9413\ : InMux
    port map (
            O => \N__38128\,
            I => \N__38121\
        );

    \I__9412\ : InMux
    port map (
            O => \N__38127\,
            I => \N__38118\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__38124\,
            I => \N__38113\
        );

    \I__9410\ : LocalMux
    port map (
            O => \N__38121\,
            I => \N__38110\
        );

    \I__9409\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38107\
        );

    \I__9408\ : InMux
    port map (
            O => \N__38117\,
            I => \N__38104\
        );

    \I__9407\ : InMux
    port map (
            O => \N__38116\,
            I => \N__38098\
        );

    \I__9406\ : Span4Mux_h
    port map (
            O => \N__38113\,
            I => \N__38093\
        );

    \I__9405\ : Span4Mux_h
    port map (
            O => \N__38110\,
            I => \N__38093\
        );

    \I__9404\ : Span4Mux_h
    port map (
            O => \N__38107\,
            I => \N__38088\
        );

    \I__9403\ : LocalMux
    port map (
            O => \N__38104\,
            I => \N__38088\
        );

    \I__9402\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38085\
        );

    \I__9401\ : InMux
    port map (
            O => \N__38102\,
            I => \N__38082\
        );

    \I__9400\ : InMux
    port map (
            O => \N__38101\,
            I => \N__38079\
        );

    \I__9399\ : LocalMux
    port map (
            O => \N__38098\,
            I => \N__38075\
        );

    \I__9398\ : Span4Mux_v
    port map (
            O => \N__38093\,
            I => \N__38072\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__38088\,
            I => \N__38069\
        );

    \I__9396\ : LocalMux
    port map (
            O => \N__38085\,
            I => \N__38066\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__38082\,
            I => \N__38061\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__38079\,
            I => \N__38061\
        );

    \I__9393\ : InMux
    port map (
            O => \N__38078\,
            I => \N__38058\
        );

    \I__9392\ : Span12Mux_h
    port map (
            O => \N__38075\,
            I => \N__38055\
        );

    \I__9391\ : Span4Mux_v
    port map (
            O => \N__38072\,
            I => \N__38052\
        );

    \I__9390\ : Span4Mux_v
    port map (
            O => \N__38069\,
            I => \N__38049\
        );

    \I__9389\ : Span4Mux_v
    port map (
            O => \N__38066\,
            I => \N__38042\
        );

    \I__9388\ : Span4Mux_s3_v
    port map (
            O => \N__38061\,
            I => \N__38042\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__38058\,
            I => \N__38042\
        );

    \I__9386\ : Span12Mux_v
    port map (
            O => \N__38055\,
            I => \N__38039\
        );

    \I__9385\ : Span4Mux_v
    port map (
            O => \N__38052\,
            I => \N__38036\
        );

    \I__9384\ : Span4Mux_h
    port map (
            O => \N__38049\,
            I => \N__38031\
        );

    \I__9383\ : Span4Mux_h
    port map (
            O => \N__38042\,
            I => \N__38031\
        );

    \I__9382\ : Odrv12
    port map (
            O => \N__38039\,
            I => port_data_c_0
        );

    \I__9381\ : Odrv4
    port map (
            O => \N__38036\,
            I => port_data_c_0
        );

    \I__9380\ : Odrv4
    port map (
            O => \N__38031\,
            I => port_data_c_0
        );

    \I__9379\ : InMux
    port map (
            O => \N__38024\,
            I => \N__38021\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__38021\,
            I => \N__38018\
        );

    \I__9377\ : Span4Mux_h
    port map (
            O => \N__38018\,
            I => \N__38015\
        );

    \I__9376\ : Odrv4
    port map (
            O => \N__38015\,
            I => \M_this_map_ram_write_data_0\
        );

    \I__9375\ : IoInMux
    port map (
            O => \N__38012\,
            I => \N__38009\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__38009\,
            I => \N__38004\
        );

    \I__9373\ : InMux
    port map (
            O => \N__38008\,
            I => \N__38001\
        );

    \I__9372\ : InMux
    port map (
            O => \N__38007\,
            I => \N__37998\
        );

    \I__9371\ : Span12Mux_s11_h
    port map (
            O => \N__38004\,
            I => \N__37993\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__38001\,
            I => \N__37990\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__37998\,
            I => \N__37987\
        );

    \I__9368\ : InMux
    port map (
            O => \N__37997\,
            I => \N__37984\
        );

    \I__9367\ : CascadeMux
    port map (
            O => \N__37996\,
            I => \N__37980\
        );

    \I__9366\ : Span12Mux_v
    port map (
            O => \N__37993\,
            I => \N__37975\
        );

    \I__9365\ : Span12Mux_v
    port map (
            O => \N__37990\,
            I => \N__37972\
        );

    \I__9364\ : Span4Mux_h
    port map (
            O => \N__37987\,
            I => \N__37969\
        );

    \I__9363\ : LocalMux
    port map (
            O => \N__37984\,
            I => \N__37966\
        );

    \I__9362\ : InMux
    port map (
            O => \N__37983\,
            I => \N__37961\
        );

    \I__9361\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37961\
        );

    \I__9360\ : InMux
    port map (
            O => \N__37979\,
            I => \N__37956\
        );

    \I__9359\ : InMux
    port map (
            O => \N__37978\,
            I => \N__37956\
        );

    \I__9358\ : Odrv12
    port map (
            O => \N__37975\,
            I => led_c_1
        );

    \I__9357\ : Odrv12
    port map (
            O => \N__37972\,
            I => led_c_1
        );

    \I__9356\ : Odrv4
    port map (
            O => \N__37969\,
            I => led_c_1
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__37966\,
            I => led_c_1
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__37961\,
            I => led_c_1
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__37956\,
            I => led_c_1
        );

    \I__9352\ : InMux
    port map (
            O => \N__37943\,
            I => \N__37940\
        );

    \I__9351\ : LocalMux
    port map (
            O => \N__37940\,
            I => \N__37935\
        );

    \I__9350\ : InMux
    port map (
            O => \N__37939\,
            I => \N__37932\
        );

    \I__9349\ : CascadeMux
    port map (
            O => \N__37938\,
            I => \N__37929\
        );

    \I__9348\ : Span4Mux_h
    port map (
            O => \N__37935\,
            I => \N__37926\
        );

    \I__9347\ : LocalMux
    port map (
            O => \N__37932\,
            I => \N__37923\
        );

    \I__9346\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37920\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__37926\,
            I => \N_466\
        );

    \I__9344\ : Odrv12
    port map (
            O => \N__37923\,
            I => \N_466\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__37920\,
            I => \N_466\
        );

    \I__9342\ : IoInMux
    port map (
            O => \N__37913\,
            I => \N__37910\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__37910\,
            I => \N__37907\
        );

    \I__9340\ : Span12Mux_s9_h
    port map (
            O => \N__37907\,
            I => \N__37904\
        );

    \I__9339\ : Span12Mux_v
    port map (
            O => \N__37904\,
            I => \N__37901\
        );

    \I__9338\ : Odrv12
    port map (
            O => \N__37901\,
            I => led_c_7
        );

    \I__9337\ : InMux
    port map (
            O => \N__37898\,
            I => \N__37895\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__37895\,
            I => \N__37892\
        );

    \I__9335\ : Span4Mux_v
    port map (
            O => \N__37892\,
            I => \N__37888\
        );

    \I__9334\ : InMux
    port map (
            O => \N__37891\,
            I => \N__37885\
        );

    \I__9333\ : Span4Mux_h
    port map (
            O => \N__37888\,
            I => \N__37880\
        );

    \I__9332\ : LocalMux
    port map (
            O => \N__37885\,
            I => \N__37880\
        );

    \I__9331\ : Span4Mux_h
    port map (
            O => \N__37880\,
            I => \N__37875\
        );

    \I__9330\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37871\
        );

    \I__9329\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37868\
        );

    \I__9328\ : Span4Mux_v
    port map (
            O => \N__37875\,
            I => \N__37865\
        );

    \I__9327\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37862\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__37871\,
            I => \N__37857\
        );

    \I__9325\ : LocalMux
    port map (
            O => \N__37868\,
            I => \N__37854\
        );

    \I__9324\ : Span4Mux_v
    port map (
            O => \N__37865\,
            I => \N__37847\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__37862\,
            I => \N__37847\
        );

    \I__9322\ : InMux
    port map (
            O => \N__37861\,
            I => \N__37844\
        );

    \I__9321\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37841\
        );

    \I__9320\ : Span4Mux_v
    port map (
            O => \N__37857\,
            I => \N__37838\
        );

    \I__9319\ : Span4Mux_v
    port map (
            O => \N__37854\,
            I => \N__37835\
        );

    \I__9318\ : InMux
    port map (
            O => \N__37853\,
            I => \N__37832\
        );

    \I__9317\ : InMux
    port map (
            O => \N__37852\,
            I => \N__37829\
        );

    \I__9316\ : Span4Mux_v
    port map (
            O => \N__37847\,
            I => \N__37826\
        );

    \I__9315\ : LocalMux
    port map (
            O => \N__37844\,
            I => \N__37823\
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__37841\,
            I => \N__37820\
        );

    \I__9313\ : Sp12to4
    port map (
            O => \N__37838\,
            I => \N__37817\
        );

    \I__9312\ : Span4Mux_h
    port map (
            O => \N__37835\,
            I => \N__37814\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__37832\,
            I => \N__37809\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__37829\,
            I => \N__37809\
        );

    \I__9309\ : Span4Mux_h
    port map (
            O => \N__37826\,
            I => \N__37804\
        );

    \I__9308\ : Span4Mux_v
    port map (
            O => \N__37823\,
            I => \N__37804\
        );

    \I__9307\ : Span12Mux_h
    port map (
            O => \N__37820\,
            I => \N__37801\
        );

    \I__9306\ : Span12Mux_h
    port map (
            O => \N__37817\,
            I => \N__37798\
        );

    \I__9305\ : Sp12to4
    port map (
            O => \N__37814\,
            I => \N__37793\
        );

    \I__9304\ : Span12Mux_h
    port map (
            O => \N__37809\,
            I => \N__37793\
        );

    \I__9303\ : Span4Mux_v
    port map (
            O => \N__37804\,
            I => \N__37790\
        );

    \I__9302\ : Span12Mux_h
    port map (
            O => \N__37801\,
            I => \N__37787\
        );

    \I__9301\ : Span12Mux_v
    port map (
            O => \N__37798\,
            I => \N__37782\
        );

    \I__9300\ : Span12Mux_h
    port map (
            O => \N__37793\,
            I => \N__37782\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__37790\,
            I => \N__37779\
        );

    \I__9298\ : Odrv12
    port map (
            O => \N__37787\,
            I => port_data_c_3
        );

    \I__9297\ : Odrv12
    port map (
            O => \N__37782\,
            I => port_data_c_3
        );

    \I__9296\ : Odrv4
    port map (
            O => \N__37779\,
            I => port_data_c_3
        );

    \I__9295\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37769\
        );

    \I__9294\ : LocalMux
    port map (
            O => \N__37769\,
            I => \M_this_map_ram_write_data_3\
        );

    \I__9293\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37763\
        );

    \I__9292\ : LocalMux
    port map (
            O => \N__37763\,
            I => \N__37760\
        );

    \I__9291\ : Span4Mux_v
    port map (
            O => \N__37760\,
            I => \N__37756\
        );

    \I__9290\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37753\
        );

    \I__9289\ : Span4Mux_h
    port map (
            O => \N__37756\,
            I => \N__37746\
        );

    \I__9288\ : LocalMux
    port map (
            O => \N__37753\,
            I => \N__37746\
        );

    \I__9287\ : InMux
    port map (
            O => \N__37752\,
            I => \N__37743\
        );

    \I__9286\ : InMux
    port map (
            O => \N__37751\,
            I => \N__37740\
        );

    \I__9285\ : Span4Mux_h
    port map (
            O => \N__37746\,
            I => \N__37736\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__37743\,
            I => \N__37731\
        );

    \I__9283\ : LocalMux
    port map (
            O => \N__37740\,
            I => \N__37728\
        );

    \I__9282\ : InMux
    port map (
            O => \N__37739\,
            I => \N__37725\
        );

    \I__9281\ : Span4Mux_v
    port map (
            O => \N__37736\,
            I => \N__37722\
        );

    \I__9280\ : InMux
    port map (
            O => \N__37735\,
            I => \N__37719\
        );

    \I__9279\ : InMux
    port map (
            O => \N__37734\,
            I => \N__37716\
        );

    \I__9278\ : Span4Mux_v
    port map (
            O => \N__37731\,
            I => \N__37712\
        );

    \I__9277\ : Span4Mux_v
    port map (
            O => \N__37728\,
            I => \N__37709\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37706\
        );

    \I__9275\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37701\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__37719\,
            I => \N__37701\
        );

    \I__9273\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37698\
        );

    \I__9272\ : InMux
    port map (
            O => \N__37715\,
            I => \N__37695\
        );

    \I__9271\ : Sp12to4
    port map (
            O => \N__37712\,
            I => \N__37689\
        );

    \I__9270\ : Sp12to4
    port map (
            O => \N__37709\,
            I => \N__37689\
        );

    \I__9269\ : Span4Mux_v
    port map (
            O => \N__37706\,
            I => \N__37686\
        );

    \I__9268\ : Span4Mux_v
    port map (
            O => \N__37701\,
            I => \N__37679\
        );

    \I__9267\ : Span4Mux_h
    port map (
            O => \N__37698\,
            I => \N__37679\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__37695\,
            I => \N__37679\
        );

    \I__9265\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37676\
        );

    \I__9264\ : Span12Mux_h
    port map (
            O => \N__37689\,
            I => \N__37671\
        );

    \I__9263\ : Sp12to4
    port map (
            O => \N__37686\,
            I => \N__37671\
        );

    \I__9262\ : IoSpan4Mux
    port map (
            O => \N__37679\,
            I => \N__37668\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__37676\,
            I => \N__37665\
        );

    \I__9260\ : Odrv12
    port map (
            O => \N__37671\,
            I => port_data_c_1
        );

    \I__9259\ : Odrv4
    port map (
            O => \N__37668\,
            I => port_data_c_1
        );

    \I__9258\ : Odrv12
    port map (
            O => \N__37665\,
            I => port_data_c_1
        );

    \I__9257\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37655\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__37655\,
            I => \M_this_map_ram_write_data_1\
        );

    \I__9255\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37646\
        );

    \I__9254\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37643\
        );

    \I__9253\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37640\
        );

    \I__9252\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37637\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__37646\,
            I => \N__37634\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__37643\,
            I => \N__37629\
        );

    \I__9249\ : LocalMux
    port map (
            O => \N__37640\,
            I => \N__37625\
        );

    \I__9248\ : LocalMux
    port map (
            O => \N__37637\,
            I => \N__37622\
        );

    \I__9247\ : Span4Mux_v
    port map (
            O => \N__37634\,
            I => \N__37619\
        );

    \I__9246\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37616\
        );

    \I__9245\ : InMux
    port map (
            O => \N__37632\,
            I => \N__37612\
        );

    \I__9244\ : Span4Mux_h
    port map (
            O => \N__37629\,
            I => \N__37608\
        );

    \I__9243\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37605\
        );

    \I__9242\ : Span4Mux_v
    port map (
            O => \N__37625\,
            I => \N__37602\
        );

    \I__9241\ : Span4Mux_v
    port map (
            O => \N__37622\,
            I => \N__37599\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__37619\,
            I => \N__37594\
        );

    \I__9239\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37594\
        );

    \I__9238\ : InMux
    port map (
            O => \N__37615\,
            I => \N__37591\
        );

    \I__9237\ : LocalMux
    port map (
            O => \N__37612\,
            I => \N__37588\
        );

    \I__9236\ : InMux
    port map (
            O => \N__37611\,
            I => \N__37585\
        );

    \I__9235\ : Span4Mux_h
    port map (
            O => \N__37608\,
            I => \N__37582\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__37605\,
            I => \N__37579\
        );

    \I__9233\ : Span4Mux_h
    port map (
            O => \N__37602\,
            I => \N__37576\
        );

    \I__9232\ : Span4Mux_h
    port map (
            O => \N__37599\,
            I => \N__37571\
        );

    \I__9231\ : Span4Mux_v
    port map (
            O => \N__37594\,
            I => \N__37571\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__37591\,
            I => \N__37568\
        );

    \I__9229\ : Span4Mux_h
    port map (
            O => \N__37588\,
            I => \N__37563\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__37585\,
            I => \N__37563\
        );

    \I__9227\ : Sp12to4
    port map (
            O => \N__37582\,
            I => \N__37560\
        );

    \I__9226\ : Span12Mux_v
    port map (
            O => \N__37579\,
            I => \N__37551\
        );

    \I__9225\ : Sp12to4
    port map (
            O => \N__37576\,
            I => \N__37551\
        );

    \I__9224\ : Sp12to4
    port map (
            O => \N__37571\,
            I => \N__37551\
        );

    \I__9223\ : Span12Mux_h
    port map (
            O => \N__37568\,
            I => \N__37551\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__37563\,
            I => \N__37548\
        );

    \I__9221\ : Span12Mux_v
    port map (
            O => \N__37560\,
            I => \N__37543\
        );

    \I__9220\ : Span12Mux_h
    port map (
            O => \N__37551\,
            I => \N__37543\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__37548\,
            I => \N__37540\
        );

    \I__9218\ : Odrv12
    port map (
            O => \N__37543\,
            I => port_data_c_2
        );

    \I__9217\ : Odrv4
    port map (
            O => \N__37540\,
            I => port_data_c_2
        );

    \I__9216\ : InMux
    port map (
            O => \N__37535\,
            I => \N__37532\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__37532\,
            I => \M_this_map_ram_write_data_2\
        );

    \I__9214\ : InMux
    port map (
            O => \N__37529\,
            I => \N__37526\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__37526\,
            I => \N__37523\
        );

    \I__9212\ : Span4Mux_v
    port map (
            O => \N__37523\,
            I => \N__37517\
        );

    \I__9211\ : InMux
    port map (
            O => \N__37522\,
            I => \N__37514\
        );

    \I__9210\ : CascadeMux
    port map (
            O => \N__37521\,
            I => \N__37511\
        );

    \I__9209\ : InMux
    port map (
            O => \N__37520\,
            I => \N__37508\
        );

    \I__9208\ : Span4Mux_v
    port map (
            O => \N__37517\,
            I => \N__37503\
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__37514\,
            I => \N__37500\
        );

    \I__9206\ : InMux
    port map (
            O => \N__37511\,
            I => \N__37496\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__37508\,
            I => \N__37493\
        );

    \I__9204\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37490\
        );

    \I__9203\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37487\
        );

    \I__9202\ : Span4Mux_v
    port map (
            O => \N__37503\,
            I => \N__37482\
        );

    \I__9201\ : Span4Mux_v
    port map (
            O => \N__37500\,
            I => \N__37482\
        );

    \I__9200\ : InMux
    port map (
            O => \N__37499\,
            I => \N__37479\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__37496\,
            I => \N__37476\
        );

    \I__9198\ : Span4Mux_v
    port map (
            O => \N__37493\,
            I => \N__37472\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__37490\,
            I => \N__37467\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__37487\,
            I => \N__37467\
        );

    \I__9195\ : Span4Mux_h
    port map (
            O => \N__37482\,
            I => \N__37463\
        );

    \I__9194\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37460\
        );

    \I__9193\ : Span4Mux_h
    port map (
            O => \N__37476\,
            I => \N__37457\
        );

    \I__9192\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37454\
        );

    \I__9191\ : Sp12to4
    port map (
            O => \N__37472\,
            I => \N__37451\
        );

    \I__9190\ : Span4Mux_v
    port map (
            O => \N__37467\,
            I => \N__37448\
        );

    \I__9189\ : InMux
    port map (
            O => \N__37466\,
            I => \N__37445\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__37463\,
            I => \N__37440\
        );

    \I__9187\ : Span4Mux_v
    port map (
            O => \N__37460\,
            I => \N__37440\
        );

    \I__9186\ : Span4Mux_v
    port map (
            O => \N__37457\,
            I => \N__37435\
        );

    \I__9185\ : LocalMux
    port map (
            O => \N__37454\,
            I => \N__37435\
        );

    \I__9184\ : Span12Mux_h
    port map (
            O => \N__37451\,
            I => \N__37432\
        );

    \I__9183\ : Sp12to4
    port map (
            O => \N__37448\,
            I => \N__37427\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37427\
        );

    \I__9181\ : Span4Mux_h
    port map (
            O => \N__37440\,
            I => \N__37422\
        );

    \I__9180\ : Span4Mux_v
    port map (
            O => \N__37435\,
            I => \N__37422\
        );

    \I__9179\ : Span12Mux_v
    port map (
            O => \N__37432\,
            I => \N__37419\
        );

    \I__9178\ : Span12Mux_h
    port map (
            O => \N__37427\,
            I => \N__37416\
        );

    \I__9177\ : Span4Mux_h
    port map (
            O => \N__37422\,
            I => \N__37413\
        );

    \I__9176\ : Odrv12
    port map (
            O => \N__37419\,
            I => port_data_c_4
        );

    \I__9175\ : Odrv12
    port map (
            O => \N__37416\,
            I => port_data_c_4
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__37413\,
            I => port_data_c_4
        );

    \I__9173\ : InMux
    port map (
            O => \N__37406\,
            I => \N__37403\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__37403\,
            I => \N__37400\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__37400\,
            I => \M_this_map_ram_write_data_4\
        );

    \I__9170\ : InMux
    port map (
            O => \N__37397\,
            I => \N__37393\
        );

    \I__9169\ : InMux
    port map (
            O => \N__37396\,
            I => \N__37390\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__37393\,
            I => \N__37385\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__37390\,
            I => \N__37382\
        );

    \I__9166\ : InMux
    port map (
            O => \N__37389\,
            I => \N__37379\
        );

    \I__9165\ : InMux
    port map (
            O => \N__37388\,
            I => \N__37376\
        );

    \I__9164\ : Span4Mux_v
    port map (
            O => \N__37385\,
            I => \N__37368\
        );

    \I__9163\ : Span4Mux_v
    port map (
            O => \N__37382\,
            I => \N__37368\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__37379\,
            I => \N__37368\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__37376\,
            I => \N__37365\
        );

    \I__9160\ : CascadeMux
    port map (
            O => \N__37375\,
            I => \N__37362\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__37368\,
            I => \N__37359\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__37365\,
            I => \N__37356\
        );

    \I__9157\ : InMux
    port map (
            O => \N__37362\,
            I => \N__37353\
        );

    \I__9156\ : Span4Mux_h
    port map (
            O => \N__37359\,
            I => \N__37344\
        );

    \I__9155\ : Span4Mux_v
    port map (
            O => \N__37356\,
            I => \N__37344\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__37353\,
            I => \N__37344\
        );

    \I__9153\ : InMux
    port map (
            O => \N__37352\,
            I => \N__37341\
        );

    \I__9152\ : InMux
    port map (
            O => \N__37351\,
            I => \N__37337\
        );

    \I__9151\ : Span4Mux_v
    port map (
            O => \N__37344\,
            I => \N__37332\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__37341\,
            I => \N__37332\
        );

    \I__9149\ : InMux
    port map (
            O => \N__37340\,
            I => \N__37328\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__37337\,
            I => \N__37325\
        );

    \I__9147\ : Span4Mux_v
    port map (
            O => \N__37332\,
            I => \N__37322\
        );

    \I__9146\ : CascadeMux
    port map (
            O => \N__37331\,
            I => \N__37319\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__37328\,
            I => \N__37316\
        );

    \I__9144\ : Span4Mux_v
    port map (
            O => \N__37325\,
            I => \N__37313\
        );

    \I__9143\ : Span4Mux_h
    port map (
            O => \N__37322\,
            I => \N__37309\
        );

    \I__9142\ : InMux
    port map (
            O => \N__37319\,
            I => \N__37306\
        );

    \I__9141\ : Span4Mux_h
    port map (
            O => \N__37316\,
            I => \N__37303\
        );

    \I__9140\ : Span4Mux_h
    port map (
            O => \N__37313\,
            I => \N__37300\
        );

    \I__9139\ : InMux
    port map (
            O => \N__37312\,
            I => \N__37297\
        );

    \I__9138\ : Span4Mux_h
    port map (
            O => \N__37309\,
            I => \N__37292\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__37306\,
            I => \N__37292\
        );

    \I__9136\ : Span4Mux_v
    port map (
            O => \N__37303\,
            I => \N__37289\
        );

    \I__9135\ : Span4Mux_h
    port map (
            O => \N__37300\,
            I => \N__37286\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__37297\,
            I => \N__37283\
        );

    \I__9133\ : Span4Mux_v
    port map (
            O => \N__37292\,
            I => \N__37280\
        );

    \I__9132\ : Sp12to4
    port map (
            O => \N__37289\,
            I => \N__37273\
        );

    \I__9131\ : Sp12to4
    port map (
            O => \N__37286\,
            I => \N__37273\
        );

    \I__9130\ : Span12Mux_s9_v
    port map (
            O => \N__37283\,
            I => \N__37273\
        );

    \I__9129\ : Span4Mux_h
    port map (
            O => \N__37280\,
            I => \N__37270\
        );

    \I__9128\ : Span12Mux_v
    port map (
            O => \N__37273\,
            I => \N__37267\
        );

    \I__9127\ : Span4Mux_h
    port map (
            O => \N__37270\,
            I => \N__37264\
        );

    \I__9126\ : Odrv12
    port map (
            O => \N__37267\,
            I => port_data_c_6
        );

    \I__9125\ : Odrv4
    port map (
            O => \N__37264\,
            I => port_data_c_6
        );

    \I__9124\ : InMux
    port map (
            O => \N__37259\,
            I => \N__37256\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__37256\,
            I => \N__37253\
        );

    \I__9122\ : Odrv4
    port map (
            O => \N__37253\,
            I => \M_this_map_ram_write_data_6\
        );

    \I__9121\ : IoInMux
    port map (
            O => \N__37250\,
            I => \N__37247\
        );

    \I__9120\ : LocalMux
    port map (
            O => \N__37247\,
            I => \N__37244\
        );

    \I__9119\ : Span4Mux_s3_v
    port map (
            O => \N__37244\,
            I => \N__37240\
        );

    \I__9118\ : CascadeMux
    port map (
            O => \N__37243\,
            I => \N__37237\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__37240\,
            I => \N__37234\
        );

    \I__9116\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37231\
        );

    \I__9115\ : Odrv4
    port map (
            O => \N__37234\,
            I => \M_this_ext_address_qZ0Z_10\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__37231\,
            I => \M_this_ext_address_qZ0Z_10\
        );

    \I__9113\ : InMux
    port map (
            O => \N__37226\,
            I => \un1_M_this_ext_address_q_cry_9\
        );

    \I__9112\ : IoInMux
    port map (
            O => \N__37223\,
            I => \N__37220\
        );

    \I__9111\ : LocalMux
    port map (
            O => \N__37220\,
            I => \N__37217\
        );

    \I__9110\ : IoSpan4Mux
    port map (
            O => \N__37217\,
            I => \N__37214\
        );

    \I__9109\ : IoSpan4Mux
    port map (
            O => \N__37214\,
            I => \N__37211\
        );

    \I__9108\ : Span4Mux_s3_v
    port map (
            O => \N__37211\,
            I => \N__37207\
        );

    \I__9107\ : CascadeMux
    port map (
            O => \N__37210\,
            I => \N__37204\
        );

    \I__9106\ : Span4Mux_v
    port map (
            O => \N__37207\,
            I => \N__37201\
        );

    \I__9105\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37198\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__37201\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__37198\,
            I => \M_this_ext_address_qZ0Z_11\
        );

    \I__9102\ : InMux
    port map (
            O => \N__37193\,
            I => \un1_M_this_ext_address_q_cry_10\
        );

    \I__9101\ : IoInMux
    port map (
            O => \N__37190\,
            I => \N__37187\
        );

    \I__9100\ : LocalMux
    port map (
            O => \N__37187\,
            I => \N__37184\
        );

    \I__9099\ : Span4Mux_s3_h
    port map (
            O => \N__37184\,
            I => \N__37181\
        );

    \I__9098\ : Span4Mux_h
    port map (
            O => \N__37181\,
            I => \N__37177\
        );

    \I__9097\ : CascadeMux
    port map (
            O => \N__37180\,
            I => \N__37174\
        );

    \I__9096\ : Span4Mux_h
    port map (
            O => \N__37177\,
            I => \N__37171\
        );

    \I__9095\ : InMux
    port map (
            O => \N__37174\,
            I => \N__37168\
        );

    \I__9094\ : Odrv4
    port map (
            O => \N__37171\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__9093\ : LocalMux
    port map (
            O => \N__37168\,
            I => \M_this_ext_address_qZ0Z_12\
        );

    \I__9092\ : InMux
    port map (
            O => \N__37163\,
            I => \un1_M_this_ext_address_q_cry_11\
        );

    \I__9091\ : IoInMux
    port map (
            O => \N__37160\,
            I => \N__37157\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__37157\,
            I => \N__37154\
        );

    \I__9089\ : Span4Mux_s2_h
    port map (
            O => \N__37154\,
            I => \N__37151\
        );

    \I__9088\ : Span4Mux_v
    port map (
            O => \N__37151\,
            I => \N__37147\
        );

    \I__9087\ : CascadeMux
    port map (
            O => \N__37150\,
            I => \N__37144\
        );

    \I__9086\ : Sp12to4
    port map (
            O => \N__37147\,
            I => \N__37141\
        );

    \I__9085\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37138\
        );

    \I__9084\ : Odrv12
    port map (
            O => \N__37141\,
            I => \M_this_ext_address_qZ0Z_13\
        );

    \I__9083\ : LocalMux
    port map (
            O => \N__37138\,
            I => \M_this_ext_address_qZ0Z_13\
        );

    \I__9082\ : InMux
    port map (
            O => \N__37133\,
            I => \un1_M_this_ext_address_q_cry_12\
        );

    \I__9081\ : IoInMux
    port map (
            O => \N__37130\,
            I => \N__37127\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__37127\,
            I => \N__37124\
        );

    \I__9079\ : IoSpan4Mux
    port map (
            O => \N__37124\,
            I => \N__37121\
        );

    \I__9078\ : Span4Mux_s2_h
    port map (
            O => \N__37121\,
            I => \N__37118\
        );

    \I__9077\ : Sp12to4
    port map (
            O => \N__37118\,
            I => \N__37114\
        );

    \I__9076\ : CascadeMux
    port map (
            O => \N__37117\,
            I => \N__37111\
        );

    \I__9075\ : Span12Mux_s11_h
    port map (
            O => \N__37114\,
            I => \N__37108\
        );

    \I__9074\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37105\
        );

    \I__9073\ : Odrv12
    port map (
            O => \N__37108\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__37105\,
            I => \M_this_ext_address_qZ0Z_14\
        );

    \I__9071\ : InMux
    port map (
            O => \N__37100\,
            I => \un1_M_this_ext_address_q_cry_13\
        );

    \I__9070\ : InMux
    port map (
            O => \N__37097\,
            I => \N__37073\
        );

    \I__9069\ : InMux
    port map (
            O => \N__37096\,
            I => \N__37073\
        );

    \I__9068\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37073\
        );

    \I__9067\ : InMux
    port map (
            O => \N__37094\,
            I => \N__37073\
        );

    \I__9066\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37064\
        );

    \I__9065\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37064\
        );

    \I__9064\ : InMux
    port map (
            O => \N__37091\,
            I => \N__37064\
        );

    \I__9063\ : InMux
    port map (
            O => \N__37090\,
            I => \N__37064\
        );

    \I__9062\ : InMux
    port map (
            O => \N__37089\,
            I => \N__37055\
        );

    \I__9061\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37055\
        );

    \I__9060\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37055\
        );

    \I__9059\ : InMux
    port map (
            O => \N__37086\,
            I => \N__37055\
        );

    \I__9058\ : InMux
    port map (
            O => \N__37085\,
            I => \N__37046\
        );

    \I__9057\ : InMux
    port map (
            O => \N__37084\,
            I => \N__37046\
        );

    \I__9056\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37046\
        );

    \I__9055\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37046\
        );

    \I__9054\ : LocalMux
    port map (
            O => \N__37073\,
            I => \N__37036\
        );

    \I__9053\ : LocalMux
    port map (
            O => \N__37064\,
            I => \N__37036\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__37055\,
            I => \N__37036\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__37046\,
            I => \N__37036\
        );

    \I__9050\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37033\
        );

    \I__9049\ : Span4Mux_v
    port map (
            O => \N__37036\,
            I => \N__37028\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__37033\,
            I => \N__37028\
        );

    \I__9047\ : Span4Mux_h
    port map (
            O => \N__37028\,
            I => \N__37025\
        );

    \I__9046\ : Odrv4
    port map (
            O => \N__37025\,
            I => \N_295\
        );

    \I__9045\ : InMux
    port map (
            O => \N__37022\,
            I => \un1_M_this_ext_address_q_cry_14\
        );

    \I__9044\ : IoInMux
    port map (
            O => \N__37019\,
            I => \N__37016\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37013\
        );

    \I__9042\ : Span4Mux_s2_h
    port map (
            O => \N__37013\,
            I => \N__37010\
        );

    \I__9041\ : Sp12to4
    port map (
            O => \N__37010\,
            I => \N__37007\
        );

    \I__9040\ : Span12Mux_v
    port map (
            O => \N__37007\,
            I => \N__37004\
        );

    \I__9039\ : Span12Mux_v
    port map (
            O => \N__37004\,
            I => \N__37000\
        );

    \I__9038\ : InMux
    port map (
            O => \N__37003\,
            I => \N__36997\
        );

    \I__9037\ : Odrv12
    port map (
            O => \N__37000\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__36997\,
            I => \M_this_ext_address_qZ0Z_15\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__36992\,
            I => \N__36988\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__36991\,
            I => \N__36985\
        );

    \I__9033\ : InMux
    port map (
            O => \N__36988\,
            I => \N__36979\
        );

    \I__9032\ : InMux
    port map (
            O => \N__36985\,
            I => \N__36979\
        );

    \I__9031\ : CascadeMux
    port map (
            O => \N__36984\,
            I => \N__36976\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__36979\,
            I => \N__36973\
        );

    \I__9029\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36970\
        );

    \I__9028\ : Odrv4
    port map (
            O => \N__36973\,
            I => \this_start_data_delay.N_231_0\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__36970\,
            I => \this_start_data_delay.N_231_0\
        );

    \I__9026\ : CascadeMux
    port map (
            O => \N__36965\,
            I => \N__36944\
        );

    \I__9025\ : CascadeMux
    port map (
            O => \N__36964\,
            I => \N__36940\
        );

    \I__9024\ : CascadeMux
    port map (
            O => \N__36963\,
            I => \N__36930\
        );

    \I__9023\ : InMux
    port map (
            O => \N__36962\,
            I => \N__36922\
        );

    \I__9022\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36922\
        );

    \I__9021\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36917\
        );

    \I__9020\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36917\
        );

    \I__9019\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36914\
        );

    \I__9018\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36911\
        );

    \I__9017\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36906\
        );

    \I__9016\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36906\
        );

    \I__9015\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36903\
        );

    \I__9014\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36898\
        );

    \I__9013\ : InMux
    port map (
            O => \N__36952\,
            I => \N__36898\
        );

    \I__9012\ : InMux
    port map (
            O => \N__36951\,
            I => \N__36895\
        );

    \I__9011\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36892\
        );

    \I__9010\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36887\
        );

    \I__9009\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36887\
        );

    \I__9008\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36884\
        );

    \I__9007\ : InMux
    port map (
            O => \N__36944\,
            I => \N__36881\
        );

    \I__9006\ : InMux
    port map (
            O => \N__36943\,
            I => \N__36878\
        );

    \I__9005\ : InMux
    port map (
            O => \N__36940\,
            I => \N__36875\
        );

    \I__9004\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36868\
        );

    \I__9003\ : InMux
    port map (
            O => \N__36938\,
            I => \N__36868\
        );

    \I__9002\ : InMux
    port map (
            O => \N__36937\,
            I => \N__36868\
        );

    \I__9001\ : InMux
    port map (
            O => \N__36936\,
            I => \N__36865\
        );

    \I__9000\ : InMux
    port map (
            O => \N__36935\,
            I => \N__36862\
        );

    \I__8999\ : InMux
    port map (
            O => \N__36934\,
            I => \N__36859\
        );

    \I__8998\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36856\
        );

    \I__8997\ : InMux
    port map (
            O => \N__36930\,
            I => \N__36851\
        );

    \I__8996\ : InMux
    port map (
            O => \N__36929\,
            I => \N__36851\
        );

    \I__8995\ : InMux
    port map (
            O => \N__36928\,
            I => \N__36846\
        );

    \I__8994\ : InMux
    port map (
            O => \N__36927\,
            I => \N__36846\
        );

    \I__8993\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36809\
        );

    \I__8992\ : LocalMux
    port map (
            O => \N__36917\,
            I => \N__36806\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__36914\,
            I => \N__36803\
        );

    \I__8990\ : LocalMux
    port map (
            O => \N__36911\,
            I => \N__36800\
        );

    \I__8989\ : LocalMux
    port map (
            O => \N__36906\,
            I => \N__36797\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__36903\,
            I => \N__36794\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__36898\,
            I => \N__36791\
        );

    \I__8986\ : LocalMux
    port map (
            O => \N__36895\,
            I => \N__36788\
        );

    \I__8985\ : LocalMux
    port map (
            O => \N__36892\,
            I => \N__36785\
        );

    \I__8984\ : LocalMux
    port map (
            O => \N__36887\,
            I => \N__36782\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__36884\,
            I => \N__36779\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__36881\,
            I => \N__36776\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__36878\,
            I => \N__36773\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36770\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__36868\,
            I => \N__36767\
        );

    \I__8978\ : LocalMux
    port map (
            O => \N__36865\,
            I => \N__36764\
        );

    \I__8977\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36761\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__36859\,
            I => \N__36758\
        );

    \I__8975\ : LocalMux
    port map (
            O => \N__36856\,
            I => \N__36755\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__36851\,
            I => \N__36752\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__36846\,
            I => \N__36749\
        );

    \I__8972\ : SRMux
    port map (
            O => \N__36845\,
            I => \N__36638\
        );

    \I__8971\ : SRMux
    port map (
            O => \N__36844\,
            I => \N__36638\
        );

    \I__8970\ : SRMux
    port map (
            O => \N__36843\,
            I => \N__36638\
        );

    \I__8969\ : SRMux
    port map (
            O => \N__36842\,
            I => \N__36638\
        );

    \I__8968\ : SRMux
    port map (
            O => \N__36841\,
            I => \N__36638\
        );

    \I__8967\ : SRMux
    port map (
            O => \N__36840\,
            I => \N__36638\
        );

    \I__8966\ : SRMux
    port map (
            O => \N__36839\,
            I => \N__36638\
        );

    \I__8965\ : SRMux
    port map (
            O => \N__36838\,
            I => \N__36638\
        );

    \I__8964\ : SRMux
    port map (
            O => \N__36837\,
            I => \N__36638\
        );

    \I__8963\ : SRMux
    port map (
            O => \N__36836\,
            I => \N__36638\
        );

    \I__8962\ : SRMux
    port map (
            O => \N__36835\,
            I => \N__36638\
        );

    \I__8961\ : SRMux
    port map (
            O => \N__36834\,
            I => \N__36638\
        );

    \I__8960\ : SRMux
    port map (
            O => \N__36833\,
            I => \N__36638\
        );

    \I__8959\ : SRMux
    port map (
            O => \N__36832\,
            I => \N__36638\
        );

    \I__8958\ : SRMux
    port map (
            O => \N__36831\,
            I => \N__36638\
        );

    \I__8957\ : SRMux
    port map (
            O => \N__36830\,
            I => \N__36638\
        );

    \I__8956\ : SRMux
    port map (
            O => \N__36829\,
            I => \N__36638\
        );

    \I__8955\ : SRMux
    port map (
            O => \N__36828\,
            I => \N__36638\
        );

    \I__8954\ : SRMux
    port map (
            O => \N__36827\,
            I => \N__36638\
        );

    \I__8953\ : SRMux
    port map (
            O => \N__36826\,
            I => \N__36638\
        );

    \I__8952\ : SRMux
    port map (
            O => \N__36825\,
            I => \N__36638\
        );

    \I__8951\ : SRMux
    port map (
            O => \N__36824\,
            I => \N__36638\
        );

    \I__8950\ : SRMux
    port map (
            O => \N__36823\,
            I => \N__36638\
        );

    \I__8949\ : SRMux
    port map (
            O => \N__36822\,
            I => \N__36638\
        );

    \I__8948\ : SRMux
    port map (
            O => \N__36821\,
            I => \N__36638\
        );

    \I__8947\ : SRMux
    port map (
            O => \N__36820\,
            I => \N__36638\
        );

    \I__8946\ : SRMux
    port map (
            O => \N__36819\,
            I => \N__36638\
        );

    \I__8945\ : SRMux
    port map (
            O => \N__36818\,
            I => \N__36638\
        );

    \I__8944\ : SRMux
    port map (
            O => \N__36817\,
            I => \N__36638\
        );

    \I__8943\ : SRMux
    port map (
            O => \N__36816\,
            I => \N__36638\
        );

    \I__8942\ : SRMux
    port map (
            O => \N__36815\,
            I => \N__36638\
        );

    \I__8941\ : SRMux
    port map (
            O => \N__36814\,
            I => \N__36638\
        );

    \I__8940\ : SRMux
    port map (
            O => \N__36813\,
            I => \N__36638\
        );

    \I__8939\ : SRMux
    port map (
            O => \N__36812\,
            I => \N__36638\
        );

    \I__8938\ : Glb2LocalMux
    port map (
            O => \N__36809\,
            I => \N__36638\
        );

    \I__8937\ : Glb2LocalMux
    port map (
            O => \N__36806\,
            I => \N__36638\
        );

    \I__8936\ : Glb2LocalMux
    port map (
            O => \N__36803\,
            I => \N__36638\
        );

    \I__8935\ : Glb2LocalMux
    port map (
            O => \N__36800\,
            I => \N__36638\
        );

    \I__8934\ : Glb2LocalMux
    port map (
            O => \N__36797\,
            I => \N__36638\
        );

    \I__8933\ : Glb2LocalMux
    port map (
            O => \N__36794\,
            I => \N__36638\
        );

    \I__8932\ : Glb2LocalMux
    port map (
            O => \N__36791\,
            I => \N__36638\
        );

    \I__8931\ : Glb2LocalMux
    port map (
            O => \N__36788\,
            I => \N__36638\
        );

    \I__8930\ : Glb2LocalMux
    port map (
            O => \N__36785\,
            I => \N__36638\
        );

    \I__8929\ : Glb2LocalMux
    port map (
            O => \N__36782\,
            I => \N__36638\
        );

    \I__8928\ : Glb2LocalMux
    port map (
            O => \N__36779\,
            I => \N__36638\
        );

    \I__8927\ : Glb2LocalMux
    port map (
            O => \N__36776\,
            I => \N__36638\
        );

    \I__8926\ : Glb2LocalMux
    port map (
            O => \N__36773\,
            I => \N__36638\
        );

    \I__8925\ : Glb2LocalMux
    port map (
            O => \N__36770\,
            I => \N__36638\
        );

    \I__8924\ : Glb2LocalMux
    port map (
            O => \N__36767\,
            I => \N__36638\
        );

    \I__8923\ : Glb2LocalMux
    port map (
            O => \N__36764\,
            I => \N__36638\
        );

    \I__8922\ : Glb2LocalMux
    port map (
            O => \N__36761\,
            I => \N__36638\
        );

    \I__8921\ : Glb2LocalMux
    port map (
            O => \N__36758\,
            I => \N__36638\
        );

    \I__8920\ : Glb2LocalMux
    port map (
            O => \N__36755\,
            I => \N__36638\
        );

    \I__8919\ : Glb2LocalMux
    port map (
            O => \N__36752\,
            I => \N__36638\
        );

    \I__8918\ : Glb2LocalMux
    port map (
            O => \N__36749\,
            I => \N__36638\
        );

    \I__8917\ : GlobalMux
    port map (
            O => \N__36638\,
            I => \N__36635\
        );

    \I__8916\ : gio2CtrlBuf
    port map (
            O => \N__36635\,
            I => \M_this_reset_cond_out_g_0\
        );

    \I__8915\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36626\
        );

    \I__8914\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36623\
        );

    \I__8913\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36618\
        );

    \I__8912\ : InMux
    port map (
            O => \N__36629\,
            I => \N__36618\
        );

    \I__8911\ : LocalMux
    port map (
            O => \N__36626\,
            I => \N__36609\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__36623\,
            I => \N__36609\
        );

    \I__8909\ : LocalMux
    port map (
            O => \N__36618\,
            I => \N__36609\
        );

    \I__8908\ : InMux
    port map (
            O => \N__36617\,
            I => \N__36604\
        );

    \I__8907\ : InMux
    port map (
            O => \N__36616\,
            I => \N__36604\
        );

    \I__8906\ : Span12Mux_h
    port map (
            O => \N__36609\,
            I => \N__36599\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__36604\,
            I => \N__36599\
        );

    \I__8904\ : Span12Mux_v
    port map (
            O => \N__36599\,
            I => \N__36596\
        );

    \I__8903\ : Odrv12
    port map (
            O => \N__36596\,
            I => \this_start_data_delay.N_227_0\
        );

    \I__8902\ : InMux
    port map (
            O => \N__36593\,
            I => \N__36588\
        );

    \I__8901\ : InMux
    port map (
            O => \N__36592\,
            I => \N__36583\
        );

    \I__8900\ : InMux
    port map (
            O => \N__36591\,
            I => \N__36583\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__36588\,
            I => \N__36580\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__36583\,
            I => \this_start_data_delay.N_242_0\
        );

    \I__8897\ : Odrv4
    port map (
            O => \N__36580\,
            I => \this_start_data_delay.N_242_0\
        );

    \I__8896\ : CascadeMux
    port map (
            O => \N__36575\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_\
        );

    \I__8895\ : CascadeMux
    port map (
            O => \N__36572\,
            I => \N__36569\
        );

    \I__8894\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36559\
        );

    \I__8893\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36556\
        );

    \I__8892\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36553\
        );

    \I__8891\ : CascadeMux
    port map (
            O => \N__36566\,
            I => \N__36547\
        );

    \I__8890\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36540\
        );

    \I__8889\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36532\
        );

    \I__8888\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36532\
        );

    \I__8887\ : InMux
    port map (
            O => \N__36562\,
            I => \N__36532\
        );

    \I__8886\ : LocalMux
    port map (
            O => \N__36559\,
            I => \N__36527\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__36556\,
            I => \N__36527\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__36553\,
            I => \N__36524\
        );

    \I__8883\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36521\
        );

    \I__8882\ : InMux
    port map (
            O => \N__36551\,
            I => \N__36518\
        );

    \I__8881\ : InMux
    port map (
            O => \N__36550\,
            I => \N__36515\
        );

    \I__8880\ : InMux
    port map (
            O => \N__36547\,
            I => \N__36512\
        );

    \I__8879\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36509\
        );

    \I__8878\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36506\
        );

    \I__8877\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36503\
        );

    \I__8876\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36499\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__36540\,
            I => \N__36495\
        );

    \I__8874\ : InMux
    port map (
            O => \N__36539\,
            I => \N__36491\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__36532\,
            I => \N__36486\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__36527\,
            I => \N__36486\
        );

    \I__8871\ : Span4Mux_v
    port map (
            O => \N__36524\,
            I => \N__36483\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__36521\,
            I => \N__36474\
        );

    \I__8869\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36474\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__36515\,
            I => \N__36474\
        );

    \I__8867\ : LocalMux
    port map (
            O => \N__36512\,
            I => \N__36474\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__36509\,
            I => \N__36469\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36469\
        );

    \I__8864\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36466\
        );

    \I__8863\ : InMux
    port map (
            O => \N__36502\,
            I => \N__36463\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__36499\,
            I => \N__36460\
        );

    \I__8861\ : InMux
    port map (
            O => \N__36498\,
            I => \N__36457\
        );

    \I__8860\ : Span4Mux_h
    port map (
            O => \N__36495\,
            I => \N__36454\
        );

    \I__8859\ : InMux
    port map (
            O => \N__36494\,
            I => \N__36451\
        );

    \I__8858\ : LocalMux
    port map (
            O => \N__36491\,
            I => \N__36448\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__36486\,
            I => \N__36439\
        );

    \I__8856\ : Span4Mux_v
    port map (
            O => \N__36483\,
            I => \N__36439\
        );

    \I__8855\ : Span4Mux_v
    port map (
            O => \N__36474\,
            I => \N__36439\
        );

    \I__8854\ : Span4Mux_v
    port map (
            O => \N__36469\,
            I => \N__36439\
        );

    \I__8853\ : Odrv4
    port map (
            O => \N__36466\,
            I => \N_220_0\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__36463\,
            I => \N_220_0\
        );

    \I__8851\ : Odrv12
    port map (
            O => \N__36460\,
            I => \N_220_0\
        );

    \I__8850\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N_220_0\
        );

    \I__8849\ : Odrv4
    port map (
            O => \N__36454\,
            I => \N_220_0\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__36451\,
            I => \N_220_0\
        );

    \I__8847\ : Odrv12
    port map (
            O => \N__36448\,
            I => \N_220_0\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__36439\,
            I => \N_220_0\
        );

    \I__8845\ : CascadeMux
    port map (
            O => \N__36422\,
            I => \N__36418\
        );

    \I__8844\ : InMux
    port map (
            O => \N__36421\,
            I => \N__36415\
        );

    \I__8843\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36410\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__36415\,
            I => \N__36407\
        );

    \I__8841\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36404\
        );

    \I__8840\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36401\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__36410\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__36407\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8837\ : LocalMux
    port map (
            O => \N__36404\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__36401\,
            I => \M_this_state_qZ0Z_10\
        );

    \I__8835\ : IoInMux
    port map (
            O => \N__36392\,
            I => \N__36389\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__36389\,
            I => \N__36386\
        );

    \I__8833\ : Span4Mux_s1_v
    port map (
            O => \N__36386\,
            I => \N__36383\
        );

    \I__8832\ : Span4Mux_v
    port map (
            O => \N__36383\,
            I => \N__36379\
        );

    \I__8831\ : InMux
    port map (
            O => \N__36382\,
            I => \N__36376\
        );

    \I__8830\ : Odrv4
    port map (
            O => \N__36379\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__36376\,
            I => \M_this_ext_address_qZ0Z_2\
        );

    \I__8828\ : InMux
    port map (
            O => \N__36371\,
            I => \un1_M_this_ext_address_q_cry_1\
        );

    \I__8827\ : IoInMux
    port map (
            O => \N__36368\,
            I => \N__36365\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36362\
        );

    \I__8825\ : Span4Mux_s3_h
    port map (
            O => \N__36362\,
            I => \N__36359\
        );

    \I__8824\ : Span4Mux_h
    port map (
            O => \N__36359\,
            I => \N__36356\
        );

    \I__8823\ : Span4Mux_v
    port map (
            O => \N__36356\,
            I => \N__36352\
        );

    \I__8822\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36349\
        );

    \I__8821\ : Odrv4
    port map (
            O => \N__36352\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__36349\,
            I => \M_this_ext_address_qZ0Z_3\
        );

    \I__8819\ : InMux
    port map (
            O => \N__36344\,
            I => \un1_M_this_ext_address_q_cry_2\
        );

    \I__8818\ : IoInMux
    port map (
            O => \N__36341\,
            I => \N__36338\
        );

    \I__8817\ : LocalMux
    port map (
            O => \N__36338\,
            I => \N__36335\
        );

    \I__8816\ : Span4Mux_s3_h
    port map (
            O => \N__36335\,
            I => \N__36332\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__36332\,
            I => \N__36329\
        );

    \I__8814\ : Span4Mux_h
    port map (
            O => \N__36329\,
            I => \N__36325\
        );

    \I__8813\ : InMux
    port map (
            O => \N__36328\,
            I => \N__36322\
        );

    \I__8812\ : Odrv4
    port map (
            O => \N__36325\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__36322\,
            I => \M_this_ext_address_qZ0Z_4\
        );

    \I__8810\ : InMux
    port map (
            O => \N__36317\,
            I => \un1_M_this_ext_address_q_cry_3\
        );

    \I__8809\ : IoInMux
    port map (
            O => \N__36314\,
            I => \N__36311\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__36311\,
            I => \N__36308\
        );

    \I__8807\ : IoSpan4Mux
    port map (
            O => \N__36308\,
            I => \N__36305\
        );

    \I__8806\ : Span4Mux_s3_h
    port map (
            O => \N__36305\,
            I => \N__36302\
        );

    \I__8805\ : Span4Mux_h
    port map (
            O => \N__36302\,
            I => \N__36298\
        );

    \I__8804\ : InMux
    port map (
            O => \N__36301\,
            I => \N__36295\
        );

    \I__8803\ : Odrv4
    port map (
            O => \N__36298\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__36295\,
            I => \M_this_ext_address_qZ0Z_5\
        );

    \I__8801\ : InMux
    port map (
            O => \N__36290\,
            I => \un1_M_this_ext_address_q_cry_4\
        );

    \I__8800\ : IoInMux
    port map (
            O => \N__36287\,
            I => \N__36284\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__36284\,
            I => \N__36281\
        );

    \I__8798\ : IoSpan4Mux
    port map (
            O => \N__36281\,
            I => \N__36278\
        );

    \I__8797\ : IoSpan4Mux
    port map (
            O => \N__36278\,
            I => \N__36275\
        );

    \I__8796\ : Span4Mux_s0_h
    port map (
            O => \N__36275\,
            I => \N__36272\
        );

    \I__8795\ : Sp12to4
    port map (
            O => \N__36272\,
            I => \N__36268\
        );

    \I__8794\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36265\
        );

    \I__8793\ : Odrv12
    port map (
            O => \N__36268\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__36265\,
            I => \M_this_ext_address_qZ0Z_6\
        );

    \I__8791\ : InMux
    port map (
            O => \N__36260\,
            I => \un1_M_this_ext_address_q_cry_5\
        );

    \I__8790\ : IoInMux
    port map (
            O => \N__36257\,
            I => \N__36254\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__36254\,
            I => \N__36251\
        );

    \I__8788\ : Span4Mux_s2_h
    port map (
            O => \N__36251\,
            I => \N__36248\
        );

    \I__8787\ : Sp12to4
    port map (
            O => \N__36248\,
            I => \N__36245\
        );

    \I__8786\ : Span12Mux_s11_v
    port map (
            O => \N__36245\,
            I => \N__36242\
        );

    \I__8785\ : Span12Mux_v
    port map (
            O => \N__36242\,
            I => \N__36238\
        );

    \I__8784\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36235\
        );

    \I__8783\ : Odrv12
    port map (
            O => \N__36238\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__36235\,
            I => \M_this_ext_address_qZ0Z_7\
        );

    \I__8781\ : InMux
    port map (
            O => \N__36230\,
            I => \un1_M_this_ext_address_q_cry_6\
        );

    \I__8780\ : IoInMux
    port map (
            O => \N__36227\,
            I => \N__36224\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36221\
        );

    \I__8778\ : IoSpan4Mux
    port map (
            O => \N__36221\,
            I => \N__36218\
        );

    \I__8777\ : Span4Mux_s3_v
    port map (
            O => \N__36218\,
            I => \N__36214\
        );

    \I__8776\ : CascadeMux
    port map (
            O => \N__36217\,
            I => \N__36211\
        );

    \I__8775\ : Span4Mux_v
    port map (
            O => \N__36214\,
            I => \N__36208\
        );

    \I__8774\ : InMux
    port map (
            O => \N__36211\,
            I => \N__36205\
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__36208\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__36205\,
            I => \M_this_ext_address_qZ0Z_8\
        );

    \I__8771\ : InMux
    port map (
            O => \N__36200\,
            I => \bfn_21_25_0_\
        );

    \I__8770\ : IoInMux
    port map (
            O => \N__36197\,
            I => \N__36194\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__36194\,
            I => \N__36191\
        );

    \I__8768\ : Span4Mux_s3_v
    port map (
            O => \N__36191\,
            I => \N__36187\
        );

    \I__8767\ : CascadeMux
    port map (
            O => \N__36190\,
            I => \N__36184\
        );

    \I__8766\ : Span4Mux_v
    port map (
            O => \N__36187\,
            I => \N__36181\
        );

    \I__8765\ : InMux
    port map (
            O => \N__36184\,
            I => \N__36178\
        );

    \I__8764\ : Odrv4
    port map (
            O => \N__36181\,
            I => \M_this_ext_address_qZ0Z_9\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__36178\,
            I => \M_this_ext_address_qZ0Z_9\
        );

    \I__8762\ : InMux
    port map (
            O => \N__36173\,
            I => \un1_M_this_ext_address_q_cry_8\
        );

    \I__8761\ : InMux
    port map (
            O => \N__36170\,
            I => \N__36167\
        );

    \I__8760\ : LocalMux
    port map (
            O => \N__36167\,
            I => \N__36162\
        );

    \I__8759\ : InMux
    port map (
            O => \N__36166\,
            I => \N__36157\
        );

    \I__8758\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36154\
        );

    \I__8757\ : Span12Mux_h
    port map (
            O => \N__36162\,
            I => \N__36151\
        );

    \I__8756\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36148\
        );

    \I__8755\ : InMux
    port map (
            O => \N__36160\,
            I => \N__36145\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__36157\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__36154\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__8752\ : Odrv12
    port map (
            O => \N__36151\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__36148\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__36145\,
            I => \M_this_state_qZ0Z_6\
        );

    \I__8749\ : InMux
    port map (
            O => \N__36134\,
            I => \N__36131\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__36131\,
            I => \N__36127\
        );

    \I__8747\ : InMux
    port map (
            O => \N__36130\,
            I => \N__36122\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__36127\,
            I => \N__36119\
        );

    \I__8745\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36114\
        );

    \I__8744\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36114\
        );

    \I__8743\ : LocalMux
    port map (
            O => \N__36122\,
            I => \N__36111\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__36119\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__36114\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8740\ : Odrv4
    port map (
            O => \N__36111\,
            I => \M_this_state_qZ0Z_5\
        );

    \I__8739\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36101\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__36101\,
            I => \N__36098\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__36098\,
            I => \N__36094\
        );

    \I__8736\ : InMux
    port map (
            O => \N__36097\,
            I => \N__36091\
        );

    \I__8735\ : Odrv4
    port map (
            O => \N__36094\,
            I => \this_start_data_delay.N_239_0\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__36091\,
            I => \this_start_data_delay.N_239_0\
        );

    \I__8733\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36080\
        );

    \I__8732\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36077\
        );

    \I__8731\ : InMux
    port map (
            O => \N__36084\,
            I => \N__36072\
        );

    \I__8730\ : InMux
    port map (
            O => \N__36083\,
            I => \N__36072\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__36080\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__36077\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8727\ : LocalMux
    port map (
            O => \N__36072\,
            I => \M_this_state_qZ0Z_3\
        );

    \I__8726\ : InMux
    port map (
            O => \N__36065\,
            I => \N__36062\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__36062\,
            I => \N__36059\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__36059\,
            I => \N__36056\
        );

    \I__8723\ : Span4Mux_h
    port map (
            O => \N__36056\,
            I => \N__36050\
        );

    \I__8722\ : InMux
    port map (
            O => \N__36055\,
            I => \N__36047\
        );

    \I__8721\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36042\
        );

    \I__8720\ : InMux
    port map (
            O => \N__36053\,
            I => \N__36042\
        );

    \I__8719\ : Odrv4
    port map (
            O => \N__36050\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8718\ : LocalMux
    port map (
            O => \N__36047\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__36042\,
            I => \M_this_state_qZ0Z_2\
        );

    \I__8716\ : CascadeMux
    port map (
            O => \N__36035\,
            I => \N__36029\
        );

    \I__8715\ : InMux
    port map (
            O => \N__36034\,
            I => \N__36024\
        );

    \I__8714\ : InMux
    port map (
            O => \N__36033\,
            I => \N__36024\
        );

    \I__8713\ : InMux
    port map (
            O => \N__36032\,
            I => \N__36021\
        );

    \I__8712\ : InMux
    port map (
            O => \N__36029\,
            I => \N__36017\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__36024\,
            I => \N__36014\
        );

    \I__8710\ : LocalMux
    port map (
            O => \N__36021\,
            I => \N__36011\
        );

    \I__8709\ : InMux
    port map (
            O => \N__36020\,
            I => \N__36008\
        );

    \I__8708\ : LocalMux
    port map (
            O => \N__36017\,
            I => \N__36002\
        );

    \I__8707\ : Span4Mux_v
    port map (
            O => \N__36014\,
            I => \N__36002\
        );

    \I__8706\ : Span12Mux_v
    port map (
            O => \N__36011\,
            I => \N__35999\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__36008\,
            I => \N__35996\
        );

    \I__8704\ : InMux
    port map (
            O => \N__36007\,
            I => \N__35993\
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__36002\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8702\ : Odrv12
    port map (
            O => \N__35999\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8701\ : Odrv4
    port map (
            O => \N__35996\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__35993\,
            I => \M_this_state_qZ0Z_1\
        );

    \I__8699\ : InMux
    port map (
            O => \N__35984\,
            I => \N__35980\
        );

    \I__8698\ : InMux
    port map (
            O => \N__35983\,
            I => \N__35977\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__35980\,
            I => \this_start_data_delay.N_420_3\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__35977\,
            I => \this_start_data_delay.N_420_3\
        );

    \I__8695\ : InMux
    port map (
            O => \N__35972\,
            I => \N__35966\
        );

    \I__8694\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35966\
        );

    \I__8693\ : LocalMux
    port map (
            O => \N__35966\,
            I => \N__35957\
        );

    \I__8692\ : InMux
    port map (
            O => \N__35965\,
            I => \N__35954\
        );

    \I__8691\ : InMux
    port map (
            O => \N__35964\,
            I => \N__35951\
        );

    \I__8690\ : InMux
    port map (
            O => \N__35963\,
            I => \N__35948\
        );

    \I__8689\ : InMux
    port map (
            O => \N__35962\,
            I => \N__35945\
        );

    \I__8688\ : InMux
    port map (
            O => \N__35961\,
            I => \N__35942\
        );

    \I__8687\ : InMux
    port map (
            O => \N__35960\,
            I => \N__35939\
        );

    \I__8686\ : Odrv4
    port map (
            O => \N__35957\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8685\ : LocalMux
    port map (
            O => \N__35954\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__35951\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8683\ : LocalMux
    port map (
            O => \N__35948\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__35945\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8681\ : LocalMux
    port map (
            O => \N__35942\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__35939\,
            I => \this_start_data_delay.N_23_1_0\
        );

    \I__8679\ : CascadeMux
    port map (
            O => \N__35924\,
            I => \this_start_data_delay.N_344_cascade_\
        );

    \I__8678\ : InMux
    port map (
            O => \N__35921\,
            I => \N__35917\
        );

    \I__8677\ : InMux
    port map (
            O => \N__35920\,
            I => \N__35914\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__35917\,
            I => \N_465\
        );

    \I__8675\ : LocalMux
    port map (
            O => \N__35914\,
            I => \N_465\
        );

    \I__8674\ : InMux
    port map (
            O => \N__35909\,
            I => \N__35906\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__35906\,
            I => \N__35901\
        );

    \I__8672\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35896\
        );

    \I__8671\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35896\
        );

    \I__8670\ : Span4Mux_h
    port map (
            O => \N__35901\,
            I => \N__35893\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35890\
        );

    \I__8668\ : Odrv4
    port map (
            O => \N__35893\,
            I => \this_start_data_delay.N_246_0\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__35890\,
            I => \this_start_data_delay.N_246_0\
        );

    \I__8666\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35882\
        );

    \I__8665\ : LocalMux
    port map (
            O => \N__35882\,
            I => \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__35879\,
            I => \N__35875\
        );

    \I__8663\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35872\
        );

    \I__8662\ : InMux
    port map (
            O => \N__35875\,
            I => \N__35869\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__35872\,
            I => \N__35864\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__35869\,
            I => \N__35864\
        );

    \I__8659\ : Span4Mux_v
    port map (
            O => \N__35864\,
            I => \N__35861\
        );

    \I__8658\ : Odrv4
    port map (
            O => \N__35861\,
            I => \M_last_q_RNIE8SF1\
        );

    \I__8657\ : IoInMux
    port map (
            O => \N__35858\,
            I => \N__35855\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__35855\,
            I => \N__35852\
        );

    \I__8655\ : Span12Mux_s8_v
    port map (
            O => \N__35852\,
            I => \N__35848\
        );

    \I__8654\ : InMux
    port map (
            O => \N__35851\,
            I => \N__35845\
        );

    \I__8653\ : Odrv12
    port map (
            O => \N__35848\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__8652\ : LocalMux
    port map (
            O => \N__35845\,
            I => \M_this_ext_address_qZ0Z_0\
        );

    \I__8651\ : IoInMux
    port map (
            O => \N__35840\,
            I => \N__35837\
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35834\
        );

    \I__8649\ : Span4Mux_s2_v
    port map (
            O => \N__35834\,
            I => \N__35831\
        );

    \I__8648\ : Span4Mux_h
    port map (
            O => \N__35831\,
            I => \N__35828\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__35828\,
            I => \N__35824\
        );

    \I__8646\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35821\
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__35824\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__35821\,
            I => \M_this_ext_address_qZ0Z_1\
        );

    \I__8643\ : InMux
    port map (
            O => \N__35816\,
            I => \un1_M_this_ext_address_q_cry_0\
        );

    \I__8642\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35796\
        );

    \I__8641\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35796\
        );

    \I__8640\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35796\
        );

    \I__8639\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35796\
        );

    \I__8638\ : InMux
    port map (
            O => \N__35809\,
            I => \N__35787\
        );

    \I__8637\ : InMux
    port map (
            O => \N__35808\,
            I => \N__35787\
        );

    \I__8636\ : InMux
    port map (
            O => \N__35807\,
            I => \N__35787\
        );

    \I__8635\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35787\
        );

    \I__8634\ : InMux
    port map (
            O => \N__35805\,
            I => \N__35778\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35772\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__35787\,
            I => \N__35772\
        );

    \I__8631\ : InMux
    port map (
            O => \N__35786\,
            I => \N__35767\
        );

    \I__8630\ : InMux
    port map (
            O => \N__35785\,
            I => \N__35767\
        );

    \I__8629\ : InMux
    port map (
            O => \N__35784\,
            I => \N__35758\
        );

    \I__8628\ : InMux
    port map (
            O => \N__35783\,
            I => \N__35758\
        );

    \I__8627\ : InMux
    port map (
            O => \N__35782\,
            I => \N__35758\
        );

    \I__8626\ : InMux
    port map (
            O => \N__35781\,
            I => \N__35758\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__35778\,
            I => \N__35755\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__35777\,
            I => \N__35752\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__35772\,
            I => \N__35745\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__35767\,
            I => \N__35745\
        );

    \I__8621\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35745\
        );

    \I__8620\ : Span4Mux_h
    port map (
            O => \N__35755\,
            I => \N__35742\
        );

    \I__8619\ : InMux
    port map (
            O => \N__35752\,
            I => \N__35739\
        );

    \I__8618\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35736\
        );

    \I__8617\ : Odrv4
    port map (
            O => \N__35742\,
            I => \N_241_0\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__35739\,
            I => \N_241_0\
        );

    \I__8615\ : Odrv4
    port map (
            O => \N__35736\,
            I => \N_241_0\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__35729\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_\
        );

    \I__8613\ : InMux
    port map (
            O => \N__35726\,
            I => \N__35723\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__35723\,
            I => \N__35720\
        );

    \I__8611\ : Span4Mux_h
    port map (
            O => \N__35720\,
            I => \N__35717\
        );

    \I__8610\ : Odrv4
    port map (
            O => \N__35717\,
            I => \this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0\
        );

    \I__8609\ : InMux
    port map (
            O => \N__35714\,
            I => \N__35707\
        );

    \I__8608\ : CascadeMux
    port map (
            O => \N__35713\,
            I => \N__35704\
        );

    \I__8607\ : InMux
    port map (
            O => \N__35712\,
            I => \N__35701\
        );

    \I__8606\ : InMux
    port map (
            O => \N__35711\,
            I => \N__35696\
        );

    \I__8605\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35696\
        );

    \I__8604\ : LocalMux
    port map (
            O => \N__35707\,
            I => \N__35692\
        );

    \I__8603\ : InMux
    port map (
            O => \N__35704\,
            I => \N__35689\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__35701\,
            I => \N__35686\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__35696\,
            I => \N__35683\
        );

    \I__8600\ : InMux
    port map (
            O => \N__35695\,
            I => \N__35680\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__35692\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__8598\ : LocalMux
    port map (
            O => \N__35689\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__8597\ : Odrv12
    port map (
            O => \N__35686\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__35683\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__35680\,
            I => \M_this_state_qZ0Z_12\
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__35669\,
            I => \N__35666\
        );

    \I__8593\ : InMux
    port map (
            O => \N__35666\,
            I => \N__35663\
        );

    \I__8592\ : LocalMux
    port map (
            O => \N__35663\,
            I => \this_start_data_delay.N_245_0\
        );

    \I__8591\ : InMux
    port map (
            O => \N__35660\,
            I => \N__35657\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35649\
        );

    \I__8589\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35638\
        );

    \I__8588\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35638\
        );

    \I__8587\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35638\
        );

    \I__8586\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35638\
        );

    \I__8585\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35638\
        );

    \I__8584\ : Odrv12
    port map (
            O => \N__35649\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__35638\,
            I => \M_this_state_qZ0Z_7\
        );

    \I__8582\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35630\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__35630\,
            I => \N__35625\
        );

    \I__8580\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35622\
        );

    \I__8579\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35617\
        );

    \I__8578\ : Span4Mux_h
    port map (
            O => \N__35625\,
            I => \N__35612\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__35622\,
            I => \N__35612\
        );

    \I__8576\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35608\
        );

    \I__8575\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35604\
        );

    \I__8574\ : LocalMux
    port map (
            O => \N__35617\,
            I => \N__35599\
        );

    \I__8573\ : Span4Mux_h
    port map (
            O => \N__35612\,
            I => \N__35599\
        );

    \I__8572\ : InMux
    port map (
            O => \N__35611\,
            I => \N__35596\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__35608\,
            I => \N__35593\
        );

    \I__8570\ : InMux
    port map (
            O => \N__35607\,
            I => \N__35590\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__35604\,
            I => \N__35585\
        );

    \I__8568\ : Span4Mux_v
    port map (
            O => \N__35599\,
            I => \N__35585\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__35596\,
            I => \N__35582\
        );

    \I__8566\ : Odrv12
    port map (
            O => \N__35593\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__35590\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__35585\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8563\ : Odrv12
    port map (
            O => \N__35582\,
            I => \M_this_state_qZ0Z_8\
        );

    \I__8562\ : InMux
    port map (
            O => \N__35573\,
            I => \N__35570\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__35570\,
            I => \N__35567\
        );

    \I__8560\ : Sp12to4
    port map (
            O => \N__35567\,
            I => \N__35564\
        );

    \I__8559\ : Span12Mux_v
    port map (
            O => \N__35564\,
            I => \N__35561\
        );

    \I__8558\ : Odrv12
    port map (
            O => \N__35561\,
            I => port_address_in_2
        );

    \I__8557\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35555\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__35555\,
            I => \N__35552\
        );

    \I__8555\ : Span4Mux_v
    port map (
            O => \N__35552\,
            I => \N__35549\
        );

    \I__8554\ : Span4Mux_h
    port map (
            O => \N__35549\,
            I => \N__35546\
        );

    \I__8553\ : Span4Mux_h
    port map (
            O => \N__35546\,
            I => \N__35543\
        );

    \I__8552\ : Odrv4
    port map (
            O => \N__35543\,
            I => port_address_in_6
        );

    \I__8551\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35536\
        );

    \I__8550\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35533\
        );

    \I__8549\ : LocalMux
    port map (
            O => \N__35536\,
            I => \N__35530\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__35533\,
            I => \N__35527\
        );

    \I__8547\ : Odrv4
    port map (
            O => \N__35530\,
            I => \this_vga_signals_M_this_state_d28_0_a2_0_1\
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__35527\,
            I => \this_vga_signals_M_this_state_d28_0_a2_0_1\
        );

    \I__8545\ : CEMux
    port map (
            O => \N__35522\,
            I => \N__35519\
        );

    \I__8544\ : LocalMux
    port map (
            O => \N__35519\,
            I => \N__35516\
        );

    \I__8543\ : Span4Mux_h
    port map (
            O => \N__35516\,
            I => \N__35513\
        );

    \I__8542\ : Span4Mux_h
    port map (
            O => \N__35513\,
            I => \N__35510\
        );

    \I__8541\ : Odrv4
    port map (
            O => \N__35510\,
            I => \N_1264_0\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__35507\,
            I => \N__35504\
        );

    \I__8539\ : InMux
    port map (
            O => \N__35504\,
            I => \N__35500\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__35503\,
            I => \N__35497\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__35500\,
            I => \N__35494\
        );

    \I__8536\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35491\
        );

    \I__8535\ : Span4Mux_h
    port map (
            O => \N__35494\,
            I => \N__35488\
        );

    \I__8534\ : LocalMux
    port map (
            O => \N__35491\,
            I => \N__35485\
        );

    \I__8533\ : Odrv4
    port map (
            O => \N__35488\,
            I => \this_start_data_delay.N_387\
        );

    \I__8532\ : Odrv12
    port map (
            O => \N__35485\,
            I => \this_start_data_delay.N_387\
        );

    \I__8531\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35477\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__35477\,
            I => \N__35473\
        );

    \I__8529\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35470\
        );

    \I__8528\ : Span4Mux_h
    port map (
            O => \N__35473\,
            I => \N__35464\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__35470\,
            I => \N__35464\
        );

    \I__8526\ : InMux
    port map (
            O => \N__35469\,
            I => \N__35461\
        );

    \I__8525\ : Span4Mux_v
    port map (
            O => \N__35464\,
            I => \N__35454\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__35461\,
            I => \N__35454\
        );

    \I__8523\ : InMux
    port map (
            O => \N__35460\,
            I => \N__35451\
        );

    \I__8522\ : InMux
    port map (
            O => \N__35459\,
            I => \N__35448\
        );

    \I__8521\ : Span4Mux_v
    port map (
            O => \N__35454\,
            I => \N__35445\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__35451\,
            I => \N__35440\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__35448\,
            I => \N__35440\
        );

    \I__8518\ : Span4Mux_v
    port map (
            O => \N__35445\,
            I => \N__35437\
        );

    \I__8517\ : Span12Mux_h
    port map (
            O => \N__35440\,
            I => \N__35434\
        );

    \I__8516\ : IoSpan4Mux
    port map (
            O => \N__35437\,
            I => \N__35431\
        );

    \I__8515\ : Odrv12
    port map (
            O => \N__35434\,
            I => port_address_in_0
        );

    \I__8514\ : Odrv4
    port map (
            O => \N__35431\,
            I => port_address_in_0
        );

    \I__8513\ : InMux
    port map (
            O => \N__35426\,
            I => \N__35421\
        );

    \I__8512\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35418\
        );

    \I__8511\ : CascadeMux
    port map (
            O => \N__35424\,
            I => \N__35414\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__35421\,
            I => \N__35410\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__35418\,
            I => \N__35407\
        );

    \I__8508\ : InMux
    port map (
            O => \N__35417\,
            I => \N__35404\
        );

    \I__8507\ : InMux
    port map (
            O => \N__35414\,
            I => \N__35401\
        );

    \I__8506\ : InMux
    port map (
            O => \N__35413\,
            I => \N__35398\
        );

    \I__8505\ : Span4Mux_v
    port map (
            O => \N__35410\,
            I => \N__35395\
        );

    \I__8504\ : Span4Mux_h
    port map (
            O => \N__35407\,
            I => \N__35386\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__35404\,
            I => \N__35386\
        );

    \I__8502\ : LocalMux
    port map (
            O => \N__35401\,
            I => \N__35386\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__35398\,
            I => \N__35386\
        );

    \I__8500\ : Sp12to4
    port map (
            O => \N__35395\,
            I => \N__35383\
        );

    \I__8499\ : Span4Mux_v
    port map (
            O => \N__35386\,
            I => \N__35380\
        );

    \I__8498\ : Span12Mux_h
    port map (
            O => \N__35383\,
            I => \N__35377\
        );

    \I__8497\ : Sp12to4
    port map (
            O => \N__35380\,
            I => \N__35374\
        );

    \I__8496\ : Odrv12
    port map (
            O => \N__35377\,
            I => port_address_in_4
        );

    \I__8495\ : Odrv12
    port map (
            O => \N__35374\,
            I => port_address_in_4
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__35369\,
            I => \this_start_data_delay.N_337_cascade_\
        );

    \I__8493\ : InMux
    port map (
            O => \N__35366\,
            I => \N__35360\
        );

    \I__8492\ : InMux
    port map (
            O => \N__35365\,
            I => \N__35355\
        );

    \I__8491\ : InMux
    port map (
            O => \N__35364\,
            I => \N__35355\
        );

    \I__8490\ : InMux
    port map (
            O => \N__35363\,
            I => \N__35352\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__35360\,
            I => \this_start_data_delay.N_386\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__35355\,
            I => \this_start_data_delay.N_386\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__35352\,
            I => \this_start_data_delay.N_386\
        );

    \I__8486\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35337\
        );

    \I__8485\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35337\
        );

    \I__8484\ : InMux
    port map (
            O => \N__35343\,
            I => \N__35331\
        );

    \I__8483\ : InMux
    port map (
            O => \N__35342\,
            I => \N__35331\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__35337\,
            I => \N__35328\
        );

    \I__8481\ : InMux
    port map (
            O => \N__35336\,
            I => \N__35325\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__35331\,
            I => \N__35322\
        );

    \I__8479\ : Odrv12
    port map (
            O => \N__35328\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__35325\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__8477\ : Odrv4
    port map (
            O => \N__35322\,
            I => \this_vga_signals.M_vcounter_q_6_repZ0Z1\
        );

    \I__8476\ : CascadeMux
    port map (
            O => \N__35315\,
            I => \N__35308\
        );

    \I__8475\ : InMux
    port map (
            O => \N__35314\,
            I => \N__35303\
        );

    \I__8474\ : InMux
    port map (
            O => \N__35313\,
            I => \N__35298\
        );

    \I__8473\ : InMux
    port map (
            O => \N__35312\,
            I => \N__35298\
        );

    \I__8472\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35295\
        );

    \I__8471\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35292\
        );

    \I__8470\ : InMux
    port map (
            O => \N__35307\,
            I => \N__35287\
        );

    \I__8469\ : InMux
    port map (
            O => \N__35306\,
            I => \N__35287\
        );

    \I__8468\ : LocalMux
    port map (
            O => \N__35303\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__35298\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__8466\ : LocalMux
    port map (
            O => \N__35295\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__35292\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__35287\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_8\
        );

    \I__8463\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35273\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35268\
        );

    \I__8461\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35264\
        );

    \I__8460\ : InMux
    port map (
            O => \N__35271\,
            I => \N__35261\
        );

    \I__8459\ : Span4Mux_h
    port map (
            O => \N__35268\,
            I => \N__35258\
        );

    \I__8458\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35254\
        );

    \I__8457\ : LocalMux
    port map (
            O => \N__35264\,
            I => \N__35246\
        );

    \I__8456\ : LocalMux
    port map (
            O => \N__35261\,
            I => \N__35246\
        );

    \I__8455\ : Span4Mux_h
    port map (
            O => \N__35258\,
            I => \N__35243\
        );

    \I__8454\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35240\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__35254\,
            I => \N__35236\
        );

    \I__8452\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35231\
        );

    \I__8451\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35231\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__35251\,
            I => \N__35227\
        );

    \I__8449\ : Span12Mux_h
    port map (
            O => \N__35246\,
            I => \N__35224\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__35243\,
            I => \N__35221\
        );

    \I__8447\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35218\
        );

    \I__8446\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35215\
        );

    \I__8445\ : Span4Mux_v
    port map (
            O => \N__35236\,
            I => \N__35210\
        );

    \I__8444\ : LocalMux
    port map (
            O => \N__35231\,
            I => \N__35210\
        );

    \I__8443\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35207\
        );

    \I__8442\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35204\
        );

    \I__8441\ : Odrv12
    port map (
            O => \N__35224\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__35221\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8439\ : Odrv12
    port map (
            O => \N__35218\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8438\ : LocalMux
    port map (
            O => \N__35215\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8437\ : Odrv4
    port map (
            O => \N__35210\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__35207\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__35204\,
            I => \this_vga_signals.M_vcounter_qZ0Z_9\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__35189\,
            I => \N__35186\
        );

    \I__8433\ : InMux
    port map (
            O => \N__35186\,
            I => \N__35177\
        );

    \I__8432\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35174\
        );

    \I__8431\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35169\
        );

    \I__8430\ : InMux
    port map (
            O => \N__35183\,
            I => \N__35169\
        );

    \I__8429\ : InMux
    port map (
            O => \N__35182\,
            I => \N__35164\
        );

    \I__8428\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35164\
        );

    \I__8427\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35161\
        );

    \I__8426\ : LocalMux
    port map (
            O => \N__35177\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__35174\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__8424\ : LocalMux
    port map (
            O => \N__35169\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__35164\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__35161\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_7\
        );

    \I__8421\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35147\
        );

    \I__8420\ : LocalMux
    port map (
            O => \N__35147\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_1\
        );

    \I__8419\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35141\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__35141\,
            I => \N__35138\
        );

    \I__8417\ : Odrv4
    port map (
            O => \N__35138\,
            I => \this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3\
        );

    \I__8416\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35132\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__35132\,
            I => \N__35127\
        );

    \I__8414\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35124\
        );

    \I__8413\ : InMux
    port map (
            O => \N__35130\,
            I => \N__35121\
        );

    \I__8412\ : Span4Mux_v
    port map (
            O => \N__35127\,
            I => \N__35117\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__35124\,
            I => \N__35112\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__35121\,
            I => \N__35112\
        );

    \I__8409\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35109\
        );

    \I__8408\ : Odrv4
    port map (
            O => \N__35117\,
            I => \this_start_data_delay.N_424\
        );

    \I__8407\ : Odrv12
    port map (
            O => \N__35112\,
            I => \this_start_data_delay.N_424\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__35109\,
            I => \this_start_data_delay.N_424\
        );

    \I__8405\ : InMux
    port map (
            O => \N__35102\,
            I => \N__35099\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__8403\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35090\
        );

    \I__8402\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35086\
        );

    \I__8401\ : InMux
    port map (
            O => \N__35096\,
            I => \N__35082\
        );

    \I__8400\ : Span4Mux_h
    port map (
            O => \N__35093\,
            I => \N__35079\
        );

    \I__8399\ : LocalMux
    port map (
            O => \N__35090\,
            I => \N__35076\
        );

    \I__8398\ : InMux
    port map (
            O => \N__35089\,
            I => \N__35073\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__35086\,
            I => \N__35069\
        );

    \I__8396\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35066\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35063\
        );

    \I__8394\ : Span4Mux_v
    port map (
            O => \N__35079\,
            I => \N__35058\
        );

    \I__8393\ : Span4Mux_h
    port map (
            O => \N__35076\,
            I => \N__35058\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__35073\,
            I => \N__35055\
        );

    \I__8391\ : InMux
    port map (
            O => \N__35072\,
            I => \N__35052\
        );

    \I__8390\ : Span12Mux_s6_v
    port map (
            O => \N__35069\,
            I => \N__35048\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__35066\,
            I => \N__35045\
        );

    \I__8388\ : Span4Mux_h
    port map (
            O => \N__35063\,
            I => \N__35042\
        );

    \I__8387\ : Span4Mux_v
    port map (
            O => \N__35058\,
            I => \N__35037\
        );

    \I__8386\ : Span4Mux_h
    port map (
            O => \N__35055\,
            I => \N__35037\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__35052\,
            I => \N__35034\
        );

    \I__8384\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35031\
        );

    \I__8383\ : Span12Mux_h
    port map (
            O => \N__35048\,
            I => \N__35028\
        );

    \I__8382\ : Span12Mux_v
    port map (
            O => \N__35045\,
            I => \N__35025\
        );

    \I__8381\ : Sp12to4
    port map (
            O => \N__35042\,
            I => \N__35022\
        );

    \I__8380\ : Span4Mux_v
    port map (
            O => \N__35037\,
            I => \N__35017\
        );

    \I__8379\ : Span4Mux_h
    port map (
            O => \N__35034\,
            I => \N__35017\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__35031\,
            I => \N__35014\
        );

    \I__8377\ : Span12Mux_v
    port map (
            O => \N__35028\,
            I => \N__35009\
        );

    \I__8376\ : Span12Mux_h
    port map (
            O => \N__35025\,
            I => \N__35009\
        );

    \I__8375\ : Span12Mux_v
    port map (
            O => \N__35022\,
            I => \N__35006\
        );

    \I__8374\ : Span4Mux_v
    port map (
            O => \N__35017\,
            I => \N__35001\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__35014\,
            I => \N__35001\
        );

    \I__8372\ : Odrv12
    port map (
            O => \N__35009\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__8371\ : Odrv12
    port map (
            O => \N__35006\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__35001\,
            I => \M_this_spr_ram_write_data_0\
        );

    \I__8369\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34990\
        );

    \I__8368\ : InMux
    port map (
            O => \N__34993\,
            I => \N__34987\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__34990\,
            I => \N__34981\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__34987\,
            I => \N__34978\
        );

    \I__8365\ : InMux
    port map (
            O => \N__34986\,
            I => \N__34975\
        );

    \I__8364\ : InMux
    port map (
            O => \N__34985\,
            I => \N__34970\
        );

    \I__8363\ : InMux
    port map (
            O => \N__34984\,
            I => \N__34967\
        );

    \I__8362\ : Span12Mux_h
    port map (
            O => \N__34981\,
            I => \N__34964\
        );

    \I__8361\ : Span4Mux_h
    port map (
            O => \N__34978\,
            I => \N__34959\
        );

    \I__8360\ : LocalMux
    port map (
            O => \N__34975\,
            I => \N__34959\
        );

    \I__8359\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34954\
        );

    \I__8358\ : InMux
    port map (
            O => \N__34973\,
            I => \N__34954\
        );

    \I__8357\ : LocalMux
    port map (
            O => \N__34970\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__34967\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8355\ : Odrv12
    port map (
            O => \N__34964\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8354\ : Odrv4
    port map (
            O => \N__34959\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__34954\,
            I => \M_this_state_qZ0Z_11\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__34943\,
            I => \this_start_data_delay.N_245_0_cascade_\
        );

    \I__8351\ : InMux
    port map (
            O => \N__34940\,
            I => \N__34937\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__34937\,
            I => \N__34934\
        );

    \I__8349\ : Odrv12
    port map (
            O => \N__34934\,
            I => un20_i_a4_0_a2_0_a2_1
        );

    \I__8348\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34927\
        );

    \I__8347\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34923\
        );

    \I__8346\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34920\
        );

    \I__8345\ : InMux
    port map (
            O => \N__34926\,
            I => \N__34917\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34913\
        );

    \I__8343\ : Span4Mux_v
    port map (
            O => \N__34920\,
            I => \N__34908\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__34917\,
            I => \N__34908\
        );

    \I__8341\ : CascadeMux
    port map (
            O => \N__34916\,
            I => \N__34904\
        );

    \I__8340\ : Span4Mux_v
    port map (
            O => \N__34913\,
            I => \N__34898\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__34908\,
            I => \N__34898\
        );

    \I__8338\ : CascadeMux
    port map (
            O => \N__34907\,
            I => \N__34895\
        );

    \I__8337\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34889\
        );

    \I__8336\ : InMux
    port map (
            O => \N__34903\,
            I => \N__34886\
        );

    \I__8335\ : Span4Mux_h
    port map (
            O => \N__34898\,
            I => \N__34883\
        );

    \I__8334\ : InMux
    port map (
            O => \N__34895\,
            I => \N__34880\
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__34894\,
            I => \N__34877\
        );

    \I__8332\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34872\
        );

    \I__8331\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34872\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__34889\,
            I => \N__34869\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__34886\,
            I => \N__34862\
        );

    \I__8328\ : Span4Mux_v
    port map (
            O => \N__34883\,
            I => \N__34862\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__34880\,
            I => \N__34862\
        );

    \I__8326\ : InMux
    port map (
            O => \N__34877\,
            I => \N__34859\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__34872\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8324\ : Odrv4
    port map (
            O => \N__34869\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__34862\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__34859\,
            I => \M_this_state_qZ0Z_13\
        );

    \I__8321\ : InMux
    port map (
            O => \N__34850\,
            I => \N__34847\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__34847\,
            I => \N__34844\
        );

    \I__8319\ : Odrv12
    port map (
            O => \N__34844\,
            I => un20_i_a4_0_a2_2
        );

    \I__8318\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34838\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__34838\,
            I => \N__34824\
        );

    \I__8316\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34819\
        );

    \I__8315\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34819\
        );

    \I__8314\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34814\
        );

    \I__8313\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34814\
        );

    \I__8312\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34805\
        );

    \I__8311\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34805\
        );

    \I__8310\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34805\
        );

    \I__8309\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34805\
        );

    \I__8308\ : InMux
    port map (
            O => \N__34829\,
            I => \N__34800\
        );

    \I__8307\ : InMux
    port map (
            O => \N__34828\,
            I => \N__34800\
        );

    \I__8306\ : InMux
    port map (
            O => \N__34827\,
            I => \N__34797\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__34824\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__34819\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__34814\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__34805\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__34800\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__34797\,
            I => \this_vga_signals.vaddress_c2\
        );

    \I__8299\ : CascadeMux
    port map (
            O => \N__34784\,
            I => \N__34781\
        );

    \I__8298\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34778\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__34778\,
            I => \this_vga_signals.N_13\
        );

    \I__8296\ : InMux
    port map (
            O => \N__34775\,
            I => \N__34772\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__34772\,
            I => \N__34768\
        );

    \I__8294\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34765\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__34768\,
            I => \N__34760\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34760\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__34760\,
            I => \N__34757\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__34757\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\
        );

    \I__8289\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34749\
        );

    \I__8288\ : CascadeMux
    port map (
            O => \N__34753\,
            I => \N__34746\
        );

    \I__8287\ : InMux
    port map (
            O => \N__34752\,
            I => \N__34742\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__34749\,
            I => \N__34739\
        );

    \I__8285\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34734\
        );

    \I__8284\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34734\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__34742\,
            I => \N__34725\
        );

    \I__8282\ : Span4Mux_h
    port map (
            O => \N__34739\,
            I => \N__34720\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34720\
        );

    \I__8280\ : InMux
    port map (
            O => \N__34733\,
            I => \N__34717\
        );

    \I__8279\ : InMux
    port map (
            O => \N__34732\,
            I => \N__34713\
        );

    \I__8278\ : InMux
    port map (
            O => \N__34731\,
            I => \N__34708\
        );

    \I__8277\ : InMux
    port map (
            O => \N__34730\,
            I => \N__34708\
        );

    \I__8276\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34703\
        );

    \I__8275\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34703\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__34725\,
            I => \N__34696\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__34720\,
            I => \N__34696\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34696\
        );

    \I__8271\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34693\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__34713\,
            I => \N__34686\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__34708\,
            I => \N__34686\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__34703\,
            I => \N__34686\
        );

    \I__8267\ : Span4Mux_h
    port map (
            O => \N__34696\,
            I => \N__34683\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__34693\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8265\ : Odrv12
    port map (
            O => \N__34686\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8264\ : Odrv4
    port map (
            O => \N__34683\,
            I => \this_vga_signals_M_vcounter_q_7\
        );

    \I__8263\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34673\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__34673\,
            I => \N__34669\
        );

    \I__8261\ : InMux
    port map (
            O => \N__34672\,
            I => \N__34666\
        );

    \I__8260\ : Span4Mux_h
    port map (
            O => \N__34669\,
            I => \N__34661\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__34666\,
            I => \N__34661\
        );

    \I__8258\ : Span4Mux_h
    port map (
            O => \N__34661\,
            I => \N__34658\
        );

    \I__8257\ : Odrv4
    port map (
            O => \N__34658\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\
        );

    \I__8256\ : CascadeMux
    port map (
            O => \N__34655\,
            I => \N__34652\
        );

    \I__8255\ : InMux
    port map (
            O => \N__34652\,
            I => \N__34644\
        );

    \I__8254\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34644\
        );

    \I__8253\ : InMux
    port map (
            O => \N__34650\,
            I => \N__34641\
        );

    \I__8252\ : InMux
    port map (
            O => \N__34649\,
            I => \N__34637\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__34644\,
            I => \N__34634\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34629\
        );

    \I__8249\ : CascadeMux
    port map (
            O => \N__34640\,
            I => \N__34623\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__34637\,
            I => \N__34617\
        );

    \I__8247\ : Span4Mux_h
    port map (
            O => \N__34634\,
            I => \N__34617\
        );

    \I__8246\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34614\
        );

    \I__8245\ : CascadeMux
    port map (
            O => \N__34632\,
            I => \N__34611\
        );

    \I__8244\ : Span4Mux_v
    port map (
            O => \N__34629\,
            I => \N__34608\
        );

    \I__8243\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34605\
        );

    \I__8242\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34600\
        );

    \I__8241\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34600\
        );

    \I__8240\ : InMux
    port map (
            O => \N__34623\,
            I => \N__34595\
        );

    \I__8239\ : InMux
    port map (
            O => \N__34622\,
            I => \N__34595\
        );

    \I__8238\ : Span4Mux_h
    port map (
            O => \N__34617\,
            I => \N__34592\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__34614\,
            I => \N__34589\
        );

    \I__8236\ : InMux
    port map (
            O => \N__34611\,
            I => \N__34586\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__34608\,
            I => \N__34577\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__34605\,
            I => \N__34577\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__34600\,
            I => \N__34577\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34577\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__34592\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__8230\ : Odrv12
    port map (
            O => \N__34589\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__34586\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__8228\ : Odrv4
    port map (
            O => \N__34577\,
            I => \this_vga_signals_M_vcounter_q_8\
        );

    \I__8227\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34565\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__34565\,
            I => \N__34561\
        );

    \I__8225\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34558\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__34561\,
            I => \N__34553\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34553\
        );

    \I__8222\ : Span4Mux_h
    port map (
            O => \N__34553\,
            I => \N__34550\
        );

    \I__8221\ : Odrv4
    port map (
            O => \N__34550\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\
        );

    \I__8220\ : InMux
    port map (
            O => \N__34547\,
            I => \N__34543\
        );

    \I__8219\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34540\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__34543\,
            I => \N__34536\
        );

    \I__8217\ : LocalMux
    port map (
            O => \N__34540\,
            I => \N__34533\
        );

    \I__8216\ : InMux
    port map (
            O => \N__34539\,
            I => \N__34530\
        );

    \I__8215\ : Span4Mux_h
    port map (
            O => \N__34536\,
            I => \N__34527\
        );

    \I__8214\ : Span4Mux_v
    port map (
            O => \N__34533\,
            I => \N__34522\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__34530\,
            I => \N__34522\
        );

    \I__8212\ : Span4Mux_h
    port map (
            O => \N__34527\,
            I => \N__34519\
        );

    \I__8211\ : Span4Mux_h
    port map (
            O => \N__34522\,
            I => \N__34516\
        );

    \I__8210\ : Odrv4
    port map (
            O => \N__34519\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__8209\ : Odrv4
    port map (
            O => \N__34516\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\
        );

    \I__8208\ : CEMux
    port map (
            O => \N__34511\,
            I => \N__34505\
        );

    \I__8207\ : CEMux
    port map (
            O => \N__34510\,
            I => \N__34502\
        );

    \I__8206\ : CEMux
    port map (
            O => \N__34509\,
            I => \N__34499\
        );

    \I__8205\ : CEMux
    port map (
            O => \N__34508\,
            I => \N__34495\
        );

    \I__8204\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34492\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__34502\,
            I => \N__34488\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__34499\,
            I => \N__34485\
        );

    \I__8201\ : CEMux
    port map (
            O => \N__34498\,
            I => \N__34481\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__34495\,
            I => \N__34476\
        );

    \I__8199\ : Span4Mux_v
    port map (
            O => \N__34492\,
            I => \N__34476\
        );

    \I__8198\ : CEMux
    port map (
            O => \N__34491\,
            I => \N__34473\
        );

    \I__8197\ : Span4Mux_v
    port map (
            O => \N__34488\,
            I => \N__34468\
        );

    \I__8196\ : Span4Mux_v
    port map (
            O => \N__34485\,
            I => \N__34468\
        );

    \I__8195\ : CEMux
    port map (
            O => \N__34484\,
            I => \N__34465\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__34481\,
            I => \N__34462\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__34476\,
            I => \N__34459\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__34473\,
            I => \N__34454\
        );

    \I__8191\ : Span4Mux_h
    port map (
            O => \N__34468\,
            I => \N__34454\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__34465\,
            I => \N__34451\
        );

    \I__8189\ : Span4Mux_h
    port map (
            O => \N__34462\,
            I => \N__34448\
        );

    \I__8188\ : Span4Mux_h
    port map (
            O => \N__34459\,
            I => \N__34445\
        );

    \I__8187\ : Span4Mux_h
    port map (
            O => \N__34454\,
            I => \N__34442\
        );

    \I__8186\ : Odrv12
    port map (
            O => \N__34451\,
            I => \this_vga_signals.N_933_0\
        );

    \I__8185\ : Odrv4
    port map (
            O => \N__34448\,
            I => \this_vga_signals.N_933_0\
        );

    \I__8184\ : Odrv4
    port map (
            O => \N__34445\,
            I => \this_vga_signals.N_933_0\
        );

    \I__8183\ : Odrv4
    port map (
            O => \N__34442\,
            I => \this_vga_signals.N_933_0\
        );

    \I__8182\ : SRMux
    port map (
            O => \N__34433\,
            I => \N__34409\
        );

    \I__8181\ : SRMux
    port map (
            O => \N__34432\,
            I => \N__34409\
        );

    \I__8180\ : SRMux
    port map (
            O => \N__34431\,
            I => \N__34409\
        );

    \I__8179\ : SRMux
    port map (
            O => \N__34430\,
            I => \N__34409\
        );

    \I__8178\ : SRMux
    port map (
            O => \N__34429\,
            I => \N__34409\
        );

    \I__8177\ : SRMux
    port map (
            O => \N__34428\,
            I => \N__34409\
        );

    \I__8176\ : SRMux
    port map (
            O => \N__34427\,
            I => \N__34409\
        );

    \I__8175\ : SRMux
    port map (
            O => \N__34426\,
            I => \N__34409\
        );

    \I__8174\ : GlobalMux
    port map (
            O => \N__34409\,
            I => \N__34406\
        );

    \I__8173\ : gio2CtrlBuf
    port map (
            O => \N__34406\,
            I => \this_vga_signals.N_1188_g\
        );

    \I__8172\ : CascadeMux
    port map (
            O => \N__34403\,
            I => \N_422_2_cascade_\
        );

    \I__8171\ : IoInMux
    port map (
            O => \N__34400\,
            I => \N__34397\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__34397\,
            I => \N__34394\
        );

    \I__8169\ : Span4Mux_s0_h
    port map (
            O => \N__34394\,
            I => \N__34391\
        );

    \I__8168\ : Span4Mux_v
    port map (
            O => \N__34391\,
            I => \N__34388\
        );

    \I__8167\ : Sp12to4
    port map (
            O => \N__34388\,
            I => \N__34385\
        );

    \I__8166\ : Span12Mux_v
    port map (
            O => \N__34385\,
            I => \N__34382\
        );

    \I__8165\ : Odrv12
    port map (
            O => \N__34382\,
            I => \N_458_i\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__34379\,
            I => \N__34376\
        );

    \I__8163\ : InMux
    port map (
            O => \N__34376\,
            I => \N__34373\
        );

    \I__8162\ : LocalMux
    port map (
            O => \N__34373\,
            I => \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6\
        );

    \I__8161\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34362\
        );

    \I__8160\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34362\
        );

    \I__8159\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34357\
        );

    \I__8158\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34357\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__34362\,
            I => \M_this_substate_qZ0\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__34357\,
            I => \M_this_substate_qZ0\
        );

    \I__8155\ : InMux
    port map (
            O => \N__34352\,
            I => \N__34345\
        );

    \I__8154\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34345\
        );

    \I__8153\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34342\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__34345\,
            I => \N__34339\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__34342\,
            I => \N__34336\
        );

    \I__8150\ : Odrv4
    port map (
            O => \N__34339\,
            I => \this_start_data_delay.N_467\
        );

    \I__8149\ : Odrv12
    port map (
            O => \N__34336\,
            I => \this_start_data_delay.N_467\
        );

    \I__8148\ : CascadeMux
    port map (
            O => \N__34331\,
            I => \this_start_data_delay.N_386_cascade_\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__34328\,
            I => \N__34322\
        );

    \I__8146\ : InMux
    port map (
            O => \N__34327\,
            I => \N__34319\
        );

    \I__8145\ : InMux
    port map (
            O => \N__34326\,
            I => \N__34312\
        );

    \I__8144\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34312\
        );

    \I__8143\ : InMux
    port map (
            O => \N__34322\,
            I => \N__34312\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__34319\,
            I => \N__34307\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__34312\,
            I => \N__34307\
        );

    \I__8140\ : Span12Mux_h
    port map (
            O => \N__34307\,
            I => \N__34304\
        );

    \I__8139\ : Odrv12
    port map (
            O => \N__34304\,
            I => port_address_in_1
        );

    \I__8138\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34292\
        );

    \I__8137\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34292\
        );

    \I__8136\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34292\
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__34292\,
            I => \this_start_data_delay.N_380\
        );

    \I__8134\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34286\
        );

    \I__8133\ : LocalMux
    port map (
            O => \N__34286\,
            I => \this_start_data_delay.N_341\
        );

    \I__8132\ : InMux
    port map (
            O => \N__34283\,
            I => \N__34279\
        );

    \I__8131\ : InMux
    port map (
            O => \N__34282\,
            I => \N__34273\
        );

    \I__8130\ : LocalMux
    port map (
            O => \N__34279\,
            I => \N__34270\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34267\
        );

    \I__8128\ : InMux
    port map (
            O => \N__34277\,
            I => \N__34264\
        );

    \I__8127\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34260\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__34273\,
            I => \N__34257\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__34270\,
            I => \N__34252\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__34267\,
            I => \N__34252\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__34264\,
            I => \N__34249\
        );

    \I__8122\ : InMux
    port map (
            O => \N__34263\,
            I => \N__34246\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__34260\,
            I => \N__34241\
        );

    \I__8120\ : Sp12to4
    port map (
            O => \N__34257\,
            I => \N__34238\
        );

    \I__8119\ : Span4Mux_v
    port map (
            O => \N__34252\,
            I => \N__34235\
        );

    \I__8118\ : Span4Mux_h
    port map (
            O => \N__34249\,
            I => \N__34232\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__34246\,
            I => \N__34229\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34226\
        );

    \I__8115\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34223\
        );

    \I__8114\ : Span12Mux_s8_h
    port map (
            O => \N__34241\,
            I => \N__34220\
        );

    \I__8113\ : Span12Mux_v
    port map (
            O => \N__34238\,
            I => \N__34217\
        );

    \I__8112\ : Sp12to4
    port map (
            O => \N__34235\,
            I => \N__34214\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__34232\,
            I => \N__34209\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__34229\,
            I => \N__34209\
        );

    \I__8109\ : LocalMux
    port map (
            O => \N__34226\,
            I => \N__34206\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__34223\,
            I => \N__34203\
        );

    \I__8107\ : Span12Mux_h
    port map (
            O => \N__34220\,
            I => \N__34200\
        );

    \I__8106\ : Span12Mux_h
    port map (
            O => \N__34217\,
            I => \N__34195\
        );

    \I__8105\ : Span12Mux_h
    port map (
            O => \N__34214\,
            I => \N__34195\
        );

    \I__8104\ : Span4Mux_v
    port map (
            O => \N__34209\,
            I => \N__34188\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__34206\,
            I => \N__34188\
        );

    \I__8102\ : Span4Mux_h
    port map (
            O => \N__34203\,
            I => \N__34188\
        );

    \I__8101\ : Odrv12
    port map (
            O => \N__34200\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__8100\ : Odrv12
    port map (
            O => \N__34195\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__8099\ : Odrv4
    port map (
            O => \N__34188\,
            I => \M_this_spr_ram_write_data_2\
        );

    \I__8098\ : CascadeMux
    port map (
            O => \N__34181\,
            I => \dma_axb0_cascade_\
        );

    \I__8097\ : InMux
    port map (
            O => \N__34178\,
            I => \N__34174\
        );

    \I__8096\ : IoInMux
    port map (
            O => \N__34177\,
            I => \N__34170\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__34174\,
            I => \N__34167\
        );

    \I__8094\ : InMux
    port map (
            O => \N__34173\,
            I => \N__34164\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__34170\,
            I => \N__34161\
        );

    \I__8092\ : Span4Mux_v
    port map (
            O => \N__34167\,
            I => \N__34158\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__34164\,
            I => \N__34155\
        );

    \I__8090\ : Span12Mux_s2_h
    port map (
            O => \N__34161\,
            I => \N__34150\
        );

    \I__8089\ : Sp12to4
    port map (
            O => \N__34158\,
            I => \N__34147\
        );

    \I__8088\ : Span4Mux_v
    port map (
            O => \N__34155\,
            I => \N__34144\
        );

    \I__8087\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34141\
        );

    \I__8086\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34138\
        );

    \I__8085\ : Span12Mux_h
    port map (
            O => \N__34150\,
            I => \N__34135\
        );

    \I__8084\ : Span12Mux_s8_h
    port map (
            O => \N__34147\,
            I => \N__34132\
        );

    \I__8083\ : Sp12to4
    port map (
            O => \N__34144\,
            I => \N__34129\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__34141\,
            I => \N__34124\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__34138\,
            I => \N__34124\
        );

    \I__8080\ : Span12Mux_v
    port map (
            O => \N__34135\,
            I => \N__34121\
        );

    \I__8079\ : Span12Mux_h
    port map (
            O => \N__34132\,
            I => \N__34116\
        );

    \I__8078\ : Span12Mux_h
    port map (
            O => \N__34129\,
            I => \N__34116\
        );

    \I__8077\ : Span4Mux_h
    port map (
            O => \N__34124\,
            I => \N__34113\
        );

    \I__8076\ : Odrv12
    port map (
            O => \N__34121\,
            I => dma_0
        );

    \I__8075\ : Odrv12
    port map (
            O => \N__34116\,
            I => dma_0
        );

    \I__8074\ : Odrv4
    port map (
            O => \N__34113\,
            I => dma_0
        );

    \I__8073\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34103\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__34103\,
            I => dma_axb3
        );

    \I__8071\ : CascadeMux
    port map (
            O => \N__34100\,
            I => \this_start_data_delay.N_345_cascade_\
        );

    \I__8070\ : InMux
    port map (
            O => \N__34097\,
            I => \N__34094\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__34094\,
            I => \N__34091\
        );

    \I__8068\ : Odrv12
    port map (
            O => \N__34091\,
            I => \this_start_data_delay.N_284_0\
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__34088\,
            I => \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__34085\,
            I => \this_start_data_delay.N_23_1_0_cascade_\
        );

    \I__8065\ : CascadeMux
    port map (
            O => \N__34082\,
            I => \this_start_data_delay.N_339_cascade_\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__34079\,
            I => \this_vga_signals.m47_0_1_cascade_\
        );

    \I__8063\ : CascadeMux
    port map (
            O => \N__34076\,
            I => \N__34070\
        );

    \I__8062\ : CascadeMux
    port map (
            O => \N__34075\,
            I => \N__34066\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__34074\,
            I => \N__34062\
        );

    \I__8060\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34057\
        );

    \I__8059\ : InMux
    port map (
            O => \N__34070\,
            I => \N__34054\
        );

    \I__8058\ : InMux
    port map (
            O => \N__34069\,
            I => \N__34049\
        );

    \I__8057\ : InMux
    port map (
            O => \N__34066\,
            I => \N__34049\
        );

    \I__8056\ : CascadeMux
    port map (
            O => \N__34065\,
            I => \N__34046\
        );

    \I__8055\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34042\
        );

    \I__8054\ : InMux
    port map (
            O => \N__34061\,
            I => \N__34038\
        );

    \I__8053\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34035\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__34057\,
            I => \N__34032\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__34054\,
            I => \N__34029\
        );

    \I__8050\ : LocalMux
    port map (
            O => \N__34049\,
            I => \N__34026\
        );

    \I__8049\ : InMux
    port map (
            O => \N__34046\,
            I => \N__34023\
        );

    \I__8048\ : InMux
    port map (
            O => \N__34045\,
            I => \N__34020\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__34042\,
            I => \N__34013\
        );

    \I__8046\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34009\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__34038\,
            I => \N__34006\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__34035\,
            I => \N__34001\
        );

    \I__8043\ : Span4Mux_v
    port map (
            O => \N__34032\,
            I => \N__34001\
        );

    \I__8042\ : Span4Mux_h
    port map (
            O => \N__34029\,
            I => \N__33992\
        );

    \I__8041\ : Span4Mux_v
    port map (
            O => \N__34026\,
            I => \N__33992\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__33992\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__33992\
        );

    \I__8038\ : InMux
    port map (
            O => \N__34019\,
            I => \N__33987\
        );

    \I__8037\ : InMux
    port map (
            O => \N__34018\,
            I => \N__33987\
        );

    \I__8036\ : CascadeMux
    port map (
            O => \N__34017\,
            I => \N__33984\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__34016\,
            I => \N__33981\
        );

    \I__8034\ : Span4Mux_v
    port map (
            O => \N__34013\,
            I => \N__33977\
        );

    \I__8033\ : InMux
    port map (
            O => \N__34012\,
            I => \N__33974\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__34009\,
            I => \N__33965\
        );

    \I__8031\ : Span4Mux_v
    port map (
            O => \N__34006\,
            I => \N__33965\
        );

    \I__8030\ : Span4Mux_h
    port map (
            O => \N__34001\,
            I => \N__33965\
        );

    \I__8029\ : Span4Mux_v
    port map (
            O => \N__33992\,
            I => \N__33965\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__33987\,
            I => \N__33962\
        );

    \I__8027\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33955\
        );

    \I__8026\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33955\
        );

    \I__8025\ : InMux
    port map (
            O => \N__33980\,
            I => \N__33955\
        );

    \I__8024\ : Odrv4
    port map (
            O => \N__33977\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__33974\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__8022\ : Odrv4
    port map (
            O => \N__33965\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__8021\ : Odrv4
    port map (
            O => \N__33962\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__33955\,
            I => \this_vga_signals_M_vcounter_q_6\
        );

    \I__8019\ : CascadeMux
    port map (
            O => \N__33944\,
            I => \N__33935\
        );

    \I__8018\ : CascadeMux
    port map (
            O => \N__33943\,
            I => \N__33932\
        );

    \I__8017\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33922\
        );

    \I__8016\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33919\
        );

    \I__8015\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33916\
        );

    \I__8014\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33913\
        );

    \I__8013\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33908\
        );

    \I__8012\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33908\
        );

    \I__8011\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33904\
        );

    \I__8010\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33898\
        );

    \I__8009\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33895\
        );

    \I__8008\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33890\
        );

    \I__8007\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33890\
        );

    \I__8006\ : CascadeMux
    port map (
            O => \N__33927\,
            I => \N__33887\
        );

    \I__8005\ : InMux
    port map (
            O => \N__33926\,
            I => \N__33884\
        );

    \I__8004\ : InMux
    port map (
            O => \N__33925\,
            I => \N__33881\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__33922\,
            I => \N__33878\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__33919\,
            I => \N__33868\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__33916\,
            I => \N__33868\
        );

    \I__8000\ : LocalMux
    port map (
            O => \N__33913\,
            I => \N__33865\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__33908\,
            I => \N__33862\
        );

    \I__7998\ : InMux
    port map (
            O => \N__33907\,
            I => \N__33859\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__33904\,
            I => \N__33856\
        );

    \I__7996\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33851\
        );

    \I__7995\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33851\
        );

    \I__7994\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33848\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33841\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33841\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__33890\,
            I => \N__33841\
        );

    \I__7990\ : InMux
    port map (
            O => \N__33887\,
            I => \N__33838\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33835\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__33881\,
            I => \N__33830\
        );

    \I__7987\ : Span4Mux_h
    port map (
            O => \N__33878\,
            I => \N__33830\
        );

    \I__7986\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33823\
        );

    \I__7985\ : InMux
    port map (
            O => \N__33876\,
            I => \N__33823\
        );

    \I__7984\ : InMux
    port map (
            O => \N__33875\,
            I => \N__33823\
        );

    \I__7983\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33818\
        );

    \I__7982\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33818\
        );

    \I__7981\ : Span4Mux_v
    port map (
            O => \N__33868\,
            I => \N__33807\
        );

    \I__7980\ : Span4Mux_v
    port map (
            O => \N__33865\,
            I => \N__33807\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__33862\,
            I => \N__33807\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__33859\,
            I => \N__33807\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__33856\,
            I => \N__33807\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__33851\,
            I => \N__33802\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__33848\,
            I => \N__33802\
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__33841\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__33838\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7972\ : Odrv4
    port map (
            O => \N__33835\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7971\ : Odrv4
    port map (
            O => \N__33830\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__33823\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__33818\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__33807\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7967\ : Odrv12
    port map (
            O => \N__33802\,
            I => \this_vga_signals.M_vcounter_qZ0Z_4\
        );

    \I__7966\ : CascadeMux
    port map (
            O => \N__33785\,
            I => \this_vga_signals.SUM_2_cascade_\
        );

    \I__7965\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33779\
        );

    \I__7964\ : LocalMux
    port map (
            O => \N__33779\,
            I => \this_vga_signals.g0_0_i_a7_1\
        );

    \I__7963\ : CascadeMux
    port map (
            O => \N__33776\,
            I => \N__33773\
        );

    \I__7962\ : InMux
    port map (
            O => \N__33773\,
            I => \N__33770\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__33770\,
            I => \N__33767\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__33767\,
            I => \N_88\
        );

    \I__7959\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33758\
        );

    \I__7958\ : InMux
    port map (
            O => \N__33763\,
            I => \N__33758\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__33758\,
            I => \N__33755\
        );

    \I__7956\ : Span12Mux_v
    port map (
            O => \N__33755\,
            I => \N__33752\
        );

    \I__7955\ : Span12Mux_h
    port map (
            O => \N__33752\,
            I => \N__33749\
        );

    \I__7954\ : Odrv12
    port map (
            O => \N__33749\,
            I => port_address_in_5
        );

    \I__7953\ : CascadeMux
    port map (
            O => \N__33746\,
            I => \N__33743\
        );

    \I__7952\ : InMux
    port map (
            O => \N__33743\,
            I => \N__33737\
        );

    \I__7951\ : InMux
    port map (
            O => \N__33742\,
            I => \N__33737\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__33737\,
            I => \N__33734\
        );

    \I__7949\ : Span4Mux_v
    port map (
            O => \N__33734\,
            I => \N__33731\
        );

    \I__7948\ : Sp12to4
    port map (
            O => \N__33731\,
            I => \N__33728\
        );

    \I__7947\ : Span12Mux_h
    port map (
            O => \N__33728\,
            I => \N__33725\
        );

    \I__7946\ : Span12Mux_v
    port map (
            O => \N__33725\,
            I => \N__33722\
        );

    \I__7945\ : Odrv12
    port map (
            O => \N__33722\,
            I => port_address_in_7
        );

    \I__7944\ : InMux
    port map (
            O => \N__33719\,
            I => \N__33713\
        );

    \I__7943\ : InMux
    port map (
            O => \N__33718\,
            I => \N__33713\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__33713\,
            I => \N__33710\
        );

    \I__7941\ : Span12Mux_v
    port map (
            O => \N__33710\,
            I => \N__33707\
        );

    \I__7940\ : Span12Mux_h
    port map (
            O => \N__33707\,
            I => \N__33704\
        );

    \I__7939\ : Odrv12
    port map (
            O => \N__33704\,
            I => port_address_in_3
        );

    \I__7938\ : CascadeMux
    port map (
            O => \N__33701\,
            I => \N__33698\
        );

    \I__7937\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33695\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__33695\,
            I => \N__33692\
        );

    \I__7935\ : Odrv4
    port map (
            O => \N__33692\,
            I => \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6\
        );

    \I__7934\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33684\
        );

    \I__7933\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33681\
        );

    \I__7932\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33678\
        );

    \I__7931\ : LocalMux
    port map (
            O => \N__33684\,
            I => \N__33673\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__33681\,
            I => \N__33673\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__33678\,
            I => \N__33670\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__33673\,
            I => \N__33667\
        );

    \I__7927\ : Span4Mux_h
    port map (
            O => \N__33670\,
            I => \N__33664\
        );

    \I__7926\ : Odrv4
    port map (
            O => \N__33667\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__33664\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\
        );

    \I__7924\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33653\
        );

    \I__7923\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33646\
        );

    \I__7922\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33646\
        );

    \I__7921\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33646\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__33653\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__33646\,
            I => \this_vga_signals.M_vcounter_q_4_repZ0Z1\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__33641\,
            I => \N__33637\
        );

    \I__7917\ : InMux
    port map (
            O => \N__33640\,
            I => \N__33632\
        );

    \I__7916\ : InMux
    port map (
            O => \N__33637\,
            I => \N__33625\
        );

    \I__7915\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33625\
        );

    \I__7914\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33625\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__33632\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__33625\,
            I => \this_vga_signals.M_vcounter_q_5_repZ0Z1\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__33620\,
            I => \N__33617\
        );

    \I__7910\ : InMux
    port map (
            O => \N__33617\,
            I => \N__33602\
        );

    \I__7909\ : InMux
    port map (
            O => \N__33616\,
            I => \N__33602\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33599\
        );

    \I__7907\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33596\
        );

    \I__7906\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33591\
        );

    \I__7905\ : InMux
    port map (
            O => \N__33612\,
            I => \N__33588\
        );

    \I__7904\ : InMux
    port map (
            O => \N__33611\,
            I => \N__33583\
        );

    \I__7903\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33583\
        );

    \I__7902\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33579\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33574\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33574\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__33602\,
            I => \N__33569\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__33599\,
            I => \N__33564\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__33596\,
            I => \N__33564\
        );

    \I__7896\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33561\
        );

    \I__7895\ : InMux
    port map (
            O => \N__33594\,
            I => \N__33558\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__33591\,
            I => \N__33555\
        );

    \I__7893\ : LocalMux
    port map (
            O => \N__33588\,
            I => \N__33550\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__33583\,
            I => \N__33550\
        );

    \I__7891\ : CascadeMux
    port map (
            O => \N__33582\,
            I => \N__33547\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__33579\,
            I => \N__33540\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__33574\,
            I => \N__33540\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__33573\,
            I => \N__33537\
        );

    \I__7887\ : CascadeMux
    port map (
            O => \N__33572\,
            I => \N__33533\
        );

    \I__7886\ : Span4Mux_h
    port map (
            O => \N__33569\,
            I => \N__33529\
        );

    \I__7885\ : Span12Mux_v
    port map (
            O => \N__33564\,
            I => \N__33524\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__33561\,
            I => \N__33524\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__33558\,
            I => \N__33517\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__33555\,
            I => \N__33517\
        );

    \I__7881\ : Span4Mux_h
    port map (
            O => \N__33550\,
            I => \N__33517\
        );

    \I__7880\ : InMux
    port map (
            O => \N__33547\,
            I => \N__33510\
        );

    \I__7879\ : InMux
    port map (
            O => \N__33546\,
            I => \N__33510\
        );

    \I__7878\ : InMux
    port map (
            O => \N__33545\,
            I => \N__33510\
        );

    \I__7877\ : Span4Mux_h
    port map (
            O => \N__33540\,
            I => \N__33507\
        );

    \I__7876\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33504\
        );

    \I__7875\ : InMux
    port map (
            O => \N__33536\,
            I => \N__33499\
        );

    \I__7874\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33499\
        );

    \I__7873\ : InMux
    port map (
            O => \N__33532\,
            I => \N__33496\
        );

    \I__7872\ : Odrv4
    port map (
            O => \N__33529\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7871\ : Odrv12
    port map (
            O => \N__33524\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7870\ : Odrv4
    port map (
            O => \N__33517\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__33510\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__33507\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__33504\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__33499\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__33496\,
            I => \this_vga_signals.vaddress_7\
        );

    \I__7864\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33467\
        );

    \I__7863\ : InMux
    port map (
            O => \N__33478\,
            I => \N__33467\
        );

    \I__7862\ : InMux
    port map (
            O => \N__33477\,
            I => \N__33460\
        );

    \I__7861\ : InMux
    port map (
            O => \N__33476\,
            I => \N__33460\
        );

    \I__7860\ : InMux
    port map (
            O => \N__33475\,
            I => \N__33460\
        );

    \I__7859\ : InMux
    port map (
            O => \N__33474\,
            I => \N__33455\
        );

    \I__7858\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33455\
        );

    \I__7857\ : InMux
    port map (
            O => \N__33472\,
            I => \N__33452\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__33467\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__33460\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__33455\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__33452\,
            I => \this_vga_signals.vaddress_6\
        );

    \I__7852\ : InMux
    port map (
            O => \N__33443\,
            I => \N__33436\
        );

    \I__7851\ : InMux
    port map (
            O => \N__33442\,
            I => \N__33429\
        );

    \I__7850\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33429\
        );

    \I__7849\ : InMux
    port map (
            O => \N__33440\,
            I => \N__33429\
        );

    \I__7848\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33426\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__33436\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__33429\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__33426\,
            I => \this_vga_signals.vaddress_5\
        );

    \I__7844\ : CascadeMux
    port map (
            O => \N__33419\,
            I => \this_vga_signals.vaddress_7_cascade_\
        );

    \I__7843\ : InMux
    port map (
            O => \N__33416\,
            I => \N__33404\
        );

    \I__7842\ : InMux
    port map (
            O => \N__33415\,
            I => \N__33399\
        );

    \I__7841\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33399\
        );

    \I__7840\ : InMux
    port map (
            O => \N__33413\,
            I => \N__33396\
        );

    \I__7839\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33393\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33390\
        );

    \I__7837\ : InMux
    port map (
            O => \N__33410\,
            I => \N__33385\
        );

    \I__7836\ : InMux
    port map (
            O => \N__33409\,
            I => \N__33385\
        );

    \I__7835\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33381\
        );

    \I__7834\ : InMux
    port map (
            O => \N__33407\,
            I => \N__33377\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__33404\,
            I => \N__33374\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__33399\,
            I => \N__33371\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__33396\,
            I => \N__33367\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__33393\,
            I => \N__33360\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__33390\,
            I => \N__33360\
        );

    \I__7828\ : LocalMux
    port map (
            O => \N__33385\,
            I => \N__33360\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33352\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__33381\,
            I => \N__33349\
        );

    \I__7825\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33346\
        );

    \I__7824\ : LocalMux
    port map (
            O => \N__33377\,
            I => \N__33343\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__33374\,
            I => \N__33338\
        );

    \I__7822\ : Span4Mux_h
    port map (
            O => \N__33371\,
            I => \N__33338\
        );

    \I__7821\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33335\
        );

    \I__7820\ : Span4Mux_v
    port map (
            O => \N__33367\,
            I => \N__33330\
        );

    \I__7819\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33330\
        );

    \I__7818\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33325\
        );

    \I__7817\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33325\
        );

    \I__7816\ : InMux
    port map (
            O => \N__33357\,
            I => \N__33320\
        );

    \I__7815\ : InMux
    port map (
            O => \N__33356\,
            I => \N__33320\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33317\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__33352\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7812\ : Odrv4
    port map (
            O => \N__33349\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__33346\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7810\ : Odrv4
    port map (
            O => \N__33343\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7809\ : Odrv4
    port map (
            O => \N__33338\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__33335\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7807\ : Odrv4
    port map (
            O => \N__33330\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__33325\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__33320\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__33317\,
            I => \this_vga_signals.SUM_2\
        );

    \I__7803\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33289\
        );

    \I__7802\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33284\
        );

    \I__7801\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33284\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33279\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33279\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__33289\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__33284\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__33279\,
            I => \this_vga_signals.if_m2_0\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__33272\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__33269\,
            I => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__33266\,
            I => \N__33262\
        );

    \I__7792\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33258\
        );

    \I__7791\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33255\
        );

    \I__7790\ : InMux
    port map (
            O => \N__33261\,
            I => \N__33250\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__33258\,
            I => \N__33245\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__33255\,
            I => \N__33245\
        );

    \I__7787\ : CascadeMux
    port map (
            O => \N__33254\,
            I => \N__33242\
        );

    \I__7786\ : CascadeMux
    port map (
            O => \N__33253\,
            I => \N__33239\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__33250\,
            I => \N__33234\
        );

    \I__7784\ : Span4Mux_v
    port map (
            O => \N__33245\,
            I => \N__33231\
        );

    \I__7783\ : InMux
    port map (
            O => \N__33242\,
            I => \N__33222\
        );

    \I__7782\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33222\
        );

    \I__7781\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33222\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33237\,
            I => \N__33222\
        );

    \I__7779\ : Span4Mux_h
    port map (
            O => \N__33234\,
            I => \N__33219\
        );

    \I__7778\ : Odrv4
    port map (
            O => \N__33231\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__33222\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__7776\ : Odrv4
    port map (
            O => \N__33219\,
            I => \this_vga_signals.mult1_un40_sum_c3_0\
        );

    \I__7775\ : CascadeMux
    port map (
            O => \N__33212\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_\
        );

    \I__7774\ : CascadeMux
    port map (
            O => \N__33209\,
            I => \N__33206\
        );

    \I__7773\ : InMux
    port map (
            O => \N__33206\,
            I => \N__33203\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__33203\,
            I => \N__33200\
        );

    \I__7771\ : Span4Mux_h
    port map (
            O => \N__33200\,
            I => \N__33197\
        );

    \I__7770\ : Odrv4
    port map (
            O => \N__33197\,
            I => \this_vga_signals.N_14\
        );

    \I__7769\ : InMux
    port map (
            O => \N__33194\,
            I => \N__33188\
        );

    \I__7768\ : InMux
    port map (
            O => \N__33193\,
            I => \N__33188\
        );

    \I__7767\ : LocalMux
    port map (
            O => \N__33188\,
            I => \this_vga_signals.g1_6\
        );

    \I__7766\ : CascadeMux
    port map (
            O => \N__33185\,
            I => \N__33179\
        );

    \I__7765\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33176\
        );

    \I__7764\ : CascadeMux
    port map (
            O => \N__33183\,
            I => \N__33173\
        );

    \I__7763\ : CascadeMux
    port map (
            O => \N__33182\,
            I => \N__33169\
        );

    \I__7762\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33165\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__33176\,
            I => \N__33162\
        );

    \I__7760\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33159\
        );

    \I__7759\ : InMux
    port map (
            O => \N__33172\,
            I => \N__33156\
        );

    \I__7758\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33153\
        );

    \I__7757\ : CascadeMux
    port map (
            O => \N__33168\,
            I => \N__33150\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33146\
        );

    \I__7755\ : Span4Mux_h
    port map (
            O => \N__33162\,
            I => \N__33141\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__33159\,
            I => \N__33141\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33138\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__33153\,
            I => \N__33135\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33150\,
            I => \N__33132\
        );

    \I__7750\ : CascadeMux
    port map (
            O => \N__33149\,
            I => \N__33128\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__33146\,
            I => \N__33109\
        );

    \I__7748\ : Span4Mux_v
    port map (
            O => \N__33141\,
            I => \N__33109\
        );

    \I__7747\ : Span4Mux_h
    port map (
            O => \N__33138\,
            I => \N__33109\
        );

    \I__7746\ : Span4Mux_v
    port map (
            O => \N__33135\,
            I => \N__33109\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33109\
        );

    \I__7744\ : CascadeMux
    port map (
            O => \N__33131\,
            I => \N__33106\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33102\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33097\
        );

    \I__7741\ : InMux
    port map (
            O => \N__33126\,
            I => \N__33097\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33125\,
            I => \N__33092\
        );

    \I__7739\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33092\
        );

    \I__7738\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33089\
        );

    \I__7737\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33084\
        );

    \I__7736\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33084\
        );

    \I__7735\ : CascadeMux
    port map (
            O => \N__33120\,
            I => \N__33080\
        );

    \I__7734\ : Span4Mux_h
    port map (
            O => \N__33109\,
            I => \N__33074\
        );

    \I__7733\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33071\
        );

    \I__7732\ : InMux
    port map (
            O => \N__33105\,
            I => \N__33068\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__33102\,
            I => \N__33065\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__33097\,
            I => \N__33062\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__33092\,
            I => \N__33059\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__33089\,
            I => \N__33054\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__33084\,
            I => \N__33054\
        );

    \I__7726\ : InMux
    port map (
            O => \N__33083\,
            I => \N__33051\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33080\,
            I => \N__33046\
        );

    \I__7724\ : InMux
    port map (
            O => \N__33079\,
            I => \N__33046\
        );

    \I__7723\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33041\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33077\,
            I => \N__33041\
        );

    \I__7721\ : Span4Mux_h
    port map (
            O => \N__33074\,
            I => \N__33038\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__33071\,
            I => \N__33029\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__33068\,
            I => \N__33029\
        );

    \I__7718\ : Span4Mux_h
    port map (
            O => \N__33065\,
            I => \N__33029\
        );

    \I__7717\ : Span4Mux_h
    port map (
            O => \N__33062\,
            I => \N__33029\
        );

    \I__7716\ : Span4Mux_v
    port map (
            O => \N__33059\,
            I => \N__33024\
        );

    \I__7715\ : Span4Mux_h
    port map (
            O => \N__33054\,
            I => \N__33024\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__33051\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__33046\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__33041\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7711\ : Odrv4
    port map (
            O => \N__33038\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7710\ : Odrv4
    port map (
            O => \N__33029\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__33024\,
            I => \this_vga_signals.M_vcounter_qZ0Z_5\
        );

    \I__7708\ : CascadeMux
    port map (
            O => \N__33011\,
            I => \this_vga_signals.N_7_1_0_3_cascade_\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33008\,
            I => \N__33005\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__33005\,
            I => \this_vga_signals.G_5_i_o2_0_1\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32997\
        );

    \I__7704\ : InMux
    port map (
            O => \N__33001\,
            I => \N__32993\
        );

    \I__7703\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32990\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__32997\,
            I => \N__32987\
        );

    \I__7701\ : InMux
    port map (
            O => \N__32996\,
            I => \N__32980\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__32993\,
            I => \N__32977\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__32990\,
            I => \N__32974\
        );

    \I__7698\ : Span4Mux_h
    port map (
            O => \N__32987\,
            I => \N__32971\
        );

    \I__7697\ : InMux
    port map (
            O => \N__32986\,
            I => \N__32964\
        );

    \I__7696\ : InMux
    port map (
            O => \N__32985\,
            I => \N__32964\
        );

    \I__7695\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32964\
        );

    \I__7694\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32961\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__32980\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7692\ : Odrv4
    port map (
            O => \N__32977\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7691\ : Odrv4
    port map (
            O => \N__32974\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__32971\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__32964\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__32961\,
            I => \this_vga_signals.vaddress_8\
        );

    \I__7687\ : InMux
    port map (
            O => \N__32948\,
            I => \N__32945\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32939\
        );

    \I__7685\ : InMux
    port map (
            O => \N__32944\,
            I => \N__32936\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__32943\,
            I => \N__32931\
        );

    \I__7683\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32926\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__32939\,
            I => \N__32923\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__32936\,
            I => \N__32920\
        );

    \I__7680\ : InMux
    port map (
            O => \N__32935\,
            I => \N__32917\
        );

    \I__7679\ : InMux
    port map (
            O => \N__32934\,
            I => \N__32914\
        );

    \I__7678\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32909\
        );

    \I__7677\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32909\
        );

    \I__7676\ : InMux
    port map (
            O => \N__32929\,
            I => \N__32906\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__32926\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7674\ : Odrv4
    port map (
            O => \N__32923\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__32920\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__32917\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__32914\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__32909\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__32906\,
            I => \this_vga_signals.vaddress_9\
        );

    \I__7668\ : InMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__7666\ : Odrv4
    port map (
            O => \N__32885\,
            I => \this_vga_signals.N_19_0_0\
        );

    \I__7665\ : InMux
    port map (
            O => \N__32882\,
            I => \N__32876\
        );

    \I__7664\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32873\
        );

    \I__7663\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32868\
        );

    \I__7662\ : InMux
    port map (
            O => \N__32879\,
            I => \N__32868\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__32876\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__7660\ : LocalMux
    port map (
            O => \N__32873\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__32868\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_6\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__32861\,
            I => \N__32857\
        );

    \I__7657\ : CascadeMux
    port map (
            O => \N__32860\,
            I => \N__32851\
        );

    \I__7656\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32846\
        );

    \I__7655\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32846\
        );

    \I__7654\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32843\
        );

    \I__7653\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32838\
        );

    \I__7652\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32838\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__32846\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__32843\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__32838\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_9\
        );

    \I__7648\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32827\
        );

    \I__7647\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32824\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__32827\,
            I => \this_vga_signals.m47_0_0\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__32824\,
            I => \this_vga_signals.m47_0_0\
        );

    \I__7644\ : InMux
    port map (
            O => \N__32819\,
            I => \N__32811\
        );

    \I__7643\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32808\
        );

    \I__7642\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32805\
        );

    \I__7641\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32802\
        );

    \I__7640\ : InMux
    port map (
            O => \N__32815\,
            I => \N__32798\
        );

    \I__7639\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32795\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__32811\,
            I => \N__32790\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__32808\,
            I => \N__32790\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32785\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__32802\,
            I => \N__32785\
        );

    \I__7634\ : InMux
    port map (
            O => \N__32801\,
            I => \N__32782\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__32798\,
            I => \N__32779\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32776\
        );

    \I__7631\ : Span12Mux_s6_v
    port map (
            O => \N__32790\,
            I => \N__32772\
        );

    \I__7630\ : Span12Mux_v
    port map (
            O => \N__32785\,
            I => \N__32769\
        );

    \I__7629\ : LocalMux
    port map (
            O => \N__32782\,
            I => \N__32766\
        );

    \I__7628\ : Span4Mux_h
    port map (
            O => \N__32779\,
            I => \N__32763\
        );

    \I__7627\ : Span12Mux_h
    port map (
            O => \N__32776\,
            I => \N__32760\
        );

    \I__7626\ : InMux
    port map (
            O => \N__32775\,
            I => \N__32757\
        );

    \I__7625\ : Span12Mux_h
    port map (
            O => \N__32772\,
            I => \N__32750\
        );

    \I__7624\ : Span12Mux_h
    port map (
            O => \N__32769\,
            I => \N__32750\
        );

    \I__7623\ : Span12Mux_h
    port map (
            O => \N__32766\,
            I => \N__32750\
        );

    \I__7622\ : Span4Mux_h
    port map (
            O => \N__32763\,
            I => \N__32747\
        );

    \I__7621\ : Span12Mux_v
    port map (
            O => \N__32760\,
            I => \N__32742\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32742\
        );

    \I__7619\ : Odrv12
    port map (
            O => \N__32750\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7618\ : Odrv4
    port map (
            O => \N__32747\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7617\ : Odrv12
    port map (
            O => \N__32742\,
            I => \M_this_spr_ram_write_data_3\
        );

    \I__7616\ : InMux
    port map (
            O => \N__32735\,
            I => \N__32732\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__32732\,
            I => \N__32729\
        );

    \I__7614\ : Span4Mux_h
    port map (
            O => \N__32729\,
            I => \N__32726\
        );

    \I__7613\ : Odrv4
    port map (
            O => \N__32726\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_1\
        );

    \I__7612\ : InMux
    port map (
            O => \N__32723\,
            I => \N__32720\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__32720\,
            I => \N__32717\
        );

    \I__7610\ : Span4Mux_v
    port map (
            O => \N__32717\,
            I => \N__32714\
        );

    \I__7609\ : Span4Mux_v
    port map (
            O => \N__32714\,
            I => \N__32711\
        );

    \I__7608\ : Span4Mux_h
    port map (
            O => \N__32711\,
            I => \N__32708\
        );

    \I__7607\ : Odrv4
    port map (
            O => \N__32708\,
            I => \M_this_map_ram_read_data_1\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__32705\,
            I => \N__32702\
        );

    \I__7605\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32698\
        );

    \I__7604\ : InMux
    port map (
            O => \N__32701\,
            I => \N__32695\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32690\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__32695\,
            I => \N__32684\
        );

    \I__7601\ : InMux
    port map (
            O => \N__32694\,
            I => \N__32681\
        );

    \I__7600\ : InMux
    port map (
            O => \N__32693\,
            I => \N__32677\
        );

    \I__7599\ : Span4Mux_h
    port map (
            O => \N__32690\,
            I => \N__32674\
        );

    \I__7598\ : InMux
    port map (
            O => \N__32689\,
            I => \N__32671\
        );

    \I__7597\ : InMux
    port map (
            O => \N__32688\,
            I => \N__32666\
        );

    \I__7596\ : InMux
    port map (
            O => \N__32687\,
            I => \N__32660\
        );

    \I__7595\ : Span4Mux_h
    port map (
            O => \N__32684\,
            I => \N__32655\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__32681\,
            I => \N__32655\
        );

    \I__7593\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32652\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__32677\,
            I => \N__32649\
        );

    \I__7591\ : Span4Mux_h
    port map (
            O => \N__32674\,
            I => \N__32644\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__32671\,
            I => \N__32644\
        );

    \I__7589\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32641\
        );

    \I__7588\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32638\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__32666\,
            I => \N__32635\
        );

    \I__7586\ : InMux
    port map (
            O => \N__32665\,
            I => \N__32632\
        );

    \I__7585\ : InMux
    port map (
            O => \N__32664\,
            I => \N__32627\
        );

    \I__7584\ : InMux
    port map (
            O => \N__32663\,
            I => \N__32627\
        );

    \I__7583\ : LocalMux
    port map (
            O => \N__32660\,
            I => \N__32620\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__32655\,
            I => \N__32620\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__32652\,
            I => \N__32620\
        );

    \I__7580\ : Span4Mux_v
    port map (
            O => \N__32649\,
            I => \N__32617\
        );

    \I__7579\ : Sp12to4
    port map (
            O => \N__32644\,
            I => \N__32612\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32612\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32603\
        );

    \I__7576\ : Span4Mux_h
    port map (
            O => \N__32635\,
            I => \N__32603\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32603\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__32627\,
            I => \N__32603\
        );

    \I__7573\ : Span4Mux_h
    port map (
            O => \N__32620\,
            I => \N__32600\
        );

    \I__7572\ : Sp12to4
    port map (
            O => \N__32617\,
            I => \N__32595\
        );

    \I__7571\ : Span12Mux_v
    port map (
            O => \N__32612\,
            I => \N__32595\
        );

    \I__7570\ : Odrv4
    port map (
            O => \N__32603\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__32600\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__7568\ : Odrv12
    port map (
            O => \N__32595\,
            I => \this_ppu.M_state_q_inv_1\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__32588\,
            I => \N__32584\
        );

    \I__7566\ : CascadeMux
    port map (
            O => \N__32587\,
            I => \N__32581\
        );

    \I__7565\ : InMux
    port map (
            O => \N__32584\,
            I => \N__32575\
        );

    \I__7564\ : InMux
    port map (
            O => \N__32581\,
            I => \N__32572\
        );

    \I__7563\ : CascadeMux
    port map (
            O => \N__32580\,
            I => \N__32569\
        );

    \I__7562\ : CascadeMux
    port map (
            O => \N__32579\,
            I => \N__32566\
        );

    \I__7561\ : CascadeMux
    port map (
            O => \N__32578\,
            I => \N__32558\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__32575\,
            I => \N__32550\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32550\
        );

    \I__7558\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32547\
        );

    \I__7557\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32544\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__32565\,
            I => \N__32541\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__32564\,
            I => \N__32538\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__32563\,
            I => \N__32532\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__32562\,
            I => \N__32529\
        );

    \I__7552\ : CascadeMux
    port map (
            O => \N__32561\,
            I => \N__32526\
        );

    \I__7551\ : InMux
    port map (
            O => \N__32558\,
            I => \N__32523\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__32557\,
            I => \N__32520\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__32556\,
            I => \N__32517\
        );

    \I__7548\ : CascadeMux
    port map (
            O => \N__32555\,
            I => \N__32514\
        );

    \I__7547\ : Span4Mux_s3_v
    port map (
            O => \N__32550\,
            I => \N__32507\
        );

    \I__7546\ : LocalMux
    port map (
            O => \N__32547\,
            I => \N__32507\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__32544\,
            I => \N__32507\
        );

    \I__7544\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32504\
        );

    \I__7543\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32501\
        );

    \I__7542\ : CascadeMux
    port map (
            O => \N__32537\,
            I => \N__32498\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__32536\,
            I => \N__32495\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__32535\,
            I => \N__32492\
        );

    \I__7539\ : InMux
    port map (
            O => \N__32532\,
            I => \N__32489\
        );

    \I__7538\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32486\
        );

    \I__7537\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32483\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__32523\,
            I => \N__32480\
        );

    \I__7535\ : InMux
    port map (
            O => \N__32520\,
            I => \N__32477\
        );

    \I__7534\ : InMux
    port map (
            O => \N__32517\,
            I => \N__32474\
        );

    \I__7533\ : InMux
    port map (
            O => \N__32514\,
            I => \N__32471\
        );

    \I__7532\ : Span4Mux_v
    port map (
            O => \N__32507\,
            I => \N__32464\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__32504\,
            I => \N__32464\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__32501\,
            I => \N__32464\
        );

    \I__7529\ : InMux
    port map (
            O => \N__32498\,
            I => \N__32461\
        );

    \I__7528\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32458\
        );

    \I__7527\ : InMux
    port map (
            O => \N__32492\,
            I => \N__32455\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__32489\,
            I => \N__32452\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__32486\,
            I => \N__32447\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__32483\,
            I => \N__32447\
        );

    \I__7523\ : Span12Mux_s7_v
    port map (
            O => \N__32480\,
            I => \N__32440\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__32477\,
            I => \N__32440\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32474\,
            I => \N__32440\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__32471\,
            I => \N__32437\
        );

    \I__7519\ : Span4Mux_v
    port map (
            O => \N__32464\,
            I => \N__32430\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32430\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__32458\,
            I => \N__32430\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__32455\,
            I => \N__32427\
        );

    \I__7515\ : Span12Mux_h
    port map (
            O => \N__32452\,
            I => \N__32424\
        );

    \I__7514\ : Span12Mux_v
    port map (
            O => \N__32447\,
            I => \N__32419\
        );

    \I__7513\ : Span12Mux_v
    port map (
            O => \N__32440\,
            I => \N__32419\
        );

    \I__7512\ : Span4Mux_v
    port map (
            O => \N__32437\,
            I => \N__32414\
        );

    \I__7511\ : Span4Mux_v
    port map (
            O => \N__32430\,
            I => \N__32414\
        );

    \I__7510\ : Span12Mux_h
    port map (
            O => \N__32427\,
            I => \N__32411\
        );

    \I__7509\ : Span12Mux_v
    port map (
            O => \N__32424\,
            I => \N__32406\
        );

    \I__7508\ : Span12Mux_h
    port map (
            O => \N__32419\,
            I => \N__32406\
        );

    \I__7507\ : Span4Mux_h
    port map (
            O => \N__32414\,
            I => \N__32403\
        );

    \I__7506\ : Odrv12
    port map (
            O => \N__32411\,
            I => \M_this_ppu_spr_addr_7\
        );

    \I__7505\ : Odrv12
    port map (
            O => \N__32406\,
            I => \M_this_ppu_spr_addr_7\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__32403\,
            I => \M_this_ppu_spr_addr_7\
        );

    \I__7503\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32393\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__32393\,
            I => \N__32389\
        );

    \I__7501\ : InMux
    port map (
            O => \N__32392\,
            I => \N__32386\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__32389\,
            I => \N__32382\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__32386\,
            I => \N__32379\
        );

    \I__7498\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32376\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__32382\,
            I => \N__32367\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__32379\,
            I => \N__32367\
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__32376\,
            I => \N__32364\
        );

    \I__7494\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32361\
        );

    \I__7493\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32357\
        );

    \I__7492\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32354\
        );

    \I__7491\ : InMux
    port map (
            O => \N__32372\,
            I => \N__32351\
        );

    \I__7490\ : Span4Mux_v
    port map (
            O => \N__32367\,
            I => \N__32346\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__32364\,
            I => \N__32346\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32343\
        );

    \I__7487\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32340\
        );

    \I__7486\ : LocalMux
    port map (
            O => \N__32357\,
            I => \N__32335\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32335\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__32351\,
            I => \N__32332\
        );

    \I__7483\ : Span4Mux_v
    port map (
            O => \N__32346\,
            I => \N__32327\
        );

    \I__7482\ : Span4Mux_h
    port map (
            O => \N__32343\,
            I => \N__32327\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__32340\,
            I => \N__32324\
        );

    \I__7480\ : Span12Mux_s10_v
    port map (
            O => \N__32335\,
            I => \N__32321\
        );

    \I__7479\ : Span12Mux_s9_v
    port map (
            O => \N__32332\,
            I => \N__32318\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__32327\,
            I => \N__32313\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__32324\,
            I => \N__32313\
        );

    \I__7476\ : Span12Mux_h
    port map (
            O => \N__32321\,
            I => \N__32308\
        );

    \I__7475\ : Span12Mux_h
    port map (
            O => \N__32318\,
            I => \N__32308\
        );

    \I__7474\ : Span4Mux_h
    port map (
            O => \N__32313\,
            I => \N__32305\
        );

    \I__7473\ : Odrv12
    port map (
            O => \N__32308\,
            I => \M_this_spr_ram_write_data_1\
        );

    \I__7472\ : Odrv4
    port map (
            O => \N__32305\,
            I => \M_this_spr_ram_write_data_1\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__32300\,
            I => \M_this_state_d_0_sqmuxa_2_cascade_\
        );

    \I__7470\ : CascadeMux
    port map (
            O => \N__32297\,
            I => \this_start_data_delay.N_233_0_cascade_\
        );

    \I__7469\ : CEMux
    port map (
            O => \N__32294\,
            I => \N__32291\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32287\
        );

    \I__7467\ : CEMux
    port map (
            O => \N__32290\,
            I => \N__32283\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__32287\,
            I => \N__32280\
        );

    \I__7465\ : CEMux
    port map (
            O => \N__32286\,
            I => \N__32277\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__32283\,
            I => \N__32270\
        );

    \I__7463\ : Span4Mux_h
    port map (
            O => \N__32280\,
            I => \N__32270\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__32277\,
            I => \N__32270\
        );

    \I__7461\ : Span4Mux_h
    port map (
            O => \N__32270\,
            I => \N__32267\
        );

    \I__7460\ : Odrv4
    port map (
            O => \N__32267\,
            I => \N_164\
        );

    \I__7459\ : InMux
    port map (
            O => \N__32264\,
            I => \N__32261\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__32261\,
            I => \N__32258\
        );

    \I__7457\ : Span4Mux_v
    port map (
            O => \N__32258\,
            I => \N__32255\
        );

    \I__7456\ : Odrv4
    port map (
            O => \N__32255\,
            I => \this_vga_signals.g1_3_0\
        );

    \I__7455\ : InMux
    port map (
            O => \N__32252\,
            I => \N__32249\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__32249\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6\
        );

    \I__7453\ : CEMux
    port map (
            O => \N__32246\,
            I => \N__32242\
        );

    \I__7452\ : CEMux
    port map (
            O => \N__32245\,
            I => \N__32239\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__32242\,
            I => \N__32236\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32233\
        );

    \I__7449\ : Span4Mux_v
    port map (
            O => \N__32236\,
            I => \N__32228\
        );

    \I__7448\ : Span4Mux_v
    port map (
            O => \N__32233\,
            I => \N__32228\
        );

    \I__7447\ : Span4Mux_h
    port map (
            O => \N__32228\,
            I => \N__32225\
        );

    \I__7446\ : Odrv4
    port map (
            O => \N__32225\,
            I => \this_spr_ram.mem_WE_6\
        );

    \I__7445\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32219\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__32219\,
            I => \N__32214\
        );

    \I__7443\ : InMux
    port map (
            O => \N__32218\,
            I => \N__32210\
        );

    \I__7442\ : InMux
    port map (
            O => \N__32217\,
            I => \N__32206\
        );

    \I__7441\ : Span4Mux_v
    port map (
            O => \N__32214\,
            I => \N__32201\
        );

    \I__7440\ : InMux
    port map (
            O => \N__32213\,
            I => \N__32198\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__32210\,
            I => \N__32195\
        );

    \I__7438\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32192\
        );

    \I__7437\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32189\
        );

    \I__7436\ : InMux
    port map (
            O => \N__32205\,
            I => \N__32186\
        );

    \I__7435\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32183\
        );

    \I__7434\ : Span4Mux_v
    port map (
            O => \N__32201\,
            I => \N__32178\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32178\
        );

    \I__7432\ : Span4Mux_h
    port map (
            O => \N__32195\,
            I => \N__32173\
        );

    \I__7431\ : LocalMux
    port map (
            O => \N__32192\,
            I => \N__32170\
        );

    \I__7430\ : Span4Mux_h
    port map (
            O => \N__32189\,
            I => \N__32167\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__32186\,
            I => \N__32164\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32183\,
            I => \N__32161\
        );

    \I__7427\ : Span4Mux_v
    port map (
            O => \N__32178\,
            I => \N__32158\
        );

    \I__7426\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32155\
        );

    \I__7425\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32152\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__32173\,
            I => \N__32147\
        );

    \I__7423\ : Span4Mux_v
    port map (
            O => \N__32170\,
            I => \N__32147\
        );

    \I__7422\ : Span4Mux_v
    port map (
            O => \N__32167\,
            I => \N__32140\
        );

    \I__7421\ : Span4Mux_h
    port map (
            O => \N__32164\,
            I => \N__32140\
        );

    \I__7420\ : Span4Mux_h
    port map (
            O => \N__32161\,
            I => \N__32140\
        );

    \I__7419\ : Sp12to4
    port map (
            O => \N__32158\,
            I => \N__32135\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__32155\,
            I => \N__32135\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__32152\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__7416\ : Odrv4
    port map (
            O => \N__32147\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__32140\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__7414\ : Odrv12
    port map (
            O => \N__32135\,
            I => \M_this_spr_address_qZ0Z_12\
        );

    \I__7413\ : InMux
    port map (
            O => \N__32126\,
            I => \N__32122\
        );

    \I__7412\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32119\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__32122\,
            I => \N__32113\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__32119\,
            I => \N__32110\
        );

    \I__7409\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32107\
        );

    \I__7408\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32104\
        );

    \I__7407\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32099\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__32113\,
            I => \N__32094\
        );

    \I__7405\ : Span4Mux_h
    port map (
            O => \N__32110\,
            I => \N__32094\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__32107\,
            I => \N__32091\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__32104\,
            I => \N__32088\
        );

    \I__7402\ : InMux
    port map (
            O => \N__32103\,
            I => \N__32085\
        );

    \I__7401\ : InMux
    port map (
            O => \N__32102\,
            I => \N__32082\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__32099\,
            I => \N__32077\
        );

    \I__7399\ : Span4Mux_v
    port map (
            O => \N__32094\,
            I => \N__32072\
        );

    \I__7398\ : Span4Mux_v
    port map (
            O => \N__32091\,
            I => \N__32072\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__32088\,
            I => \N__32067\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__32085\,
            I => \N__32067\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__32082\,
            I => \N__32064\
        );

    \I__7394\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32061\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32058\
        );

    \I__7392\ : Span4Mux_v
    port map (
            O => \N__32077\,
            I => \N__32055\
        );

    \I__7391\ : Span4Mux_h
    port map (
            O => \N__32072\,
            I => \N__32048\
        );

    \I__7390\ : Span4Mux_v
    port map (
            O => \N__32067\,
            I => \N__32048\
        );

    \I__7389\ : Span4Mux_v
    port map (
            O => \N__32064\,
            I => \N__32048\
        );

    \I__7388\ : LocalMux
    port map (
            O => \N__32061\,
            I => \N__32045\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__32058\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__7386\ : Odrv4
    port map (
            O => \N__32055\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__7385\ : Odrv4
    port map (
            O => \N__32048\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__7384\ : Odrv4
    port map (
            O => \N__32045\,
            I => \M_this_spr_address_qZ0Z_11\
        );

    \I__7383\ : CascadeMux
    port map (
            O => \N__32036\,
            I => \N__32033\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__32032\,
            I => \N__32024\
        );

    \I__7380\ : CascadeMux
    port map (
            O => \N__32031\,
            I => \N__32021\
        );

    \I__7379\ : CascadeMux
    port map (
            O => \N__32030\,
            I => \N__32018\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32013\
        );

    \I__7377\ : InMux
    port map (
            O => \N__32024\,
            I => \N__32010\
        );

    \I__7376\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32007\
        );

    \I__7375\ : InMux
    port map (
            O => \N__32018\,
            I => \N__32004\
        );

    \I__7374\ : CascadeMux
    port map (
            O => \N__32017\,
            I => \N__32001\
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__32016\,
            I => \N__31997\
        );

    \I__7372\ : Span4Mux_v
    port map (
            O => \N__32013\,
            I => \N__31991\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__32010\,
            I => \N__31991\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32007\,
            I => \N__31988\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31985\
        );

    \I__7368\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31982\
        );

    \I__7367\ : InMux
    port map (
            O => \N__32000\,
            I => \N__31979\
        );

    \I__7366\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31976\
        );

    \I__7365\ : CascadeMux
    port map (
            O => \N__31996\,
            I => \N__31973\
        );

    \I__7364\ : Span4Mux_h
    port map (
            O => \N__31991\,
            I => \N__31969\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__31988\,
            I => \N__31966\
        );

    \I__7362\ : Span4Mux_v
    port map (
            O => \N__31985\,
            I => \N__31963\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__31982\,
            I => \N__31960\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31957\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__31976\,
            I => \N__31954\
        );

    \I__7358\ : InMux
    port map (
            O => \N__31973\,
            I => \N__31951\
        );

    \I__7357\ : InMux
    port map (
            O => \N__31972\,
            I => \N__31948\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__31969\,
            I => \N__31941\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__31966\,
            I => \N__31941\
        );

    \I__7354\ : Span4Mux_h
    port map (
            O => \N__31963\,
            I => \N__31941\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__31960\,
            I => \N__31938\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__31957\,
            I => \N__31935\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__31954\,
            I => \N__31930\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31930\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__31948\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__7348\ : Odrv4
    port map (
            O => \N__31941\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__7347\ : Odrv4
    port map (
            O => \N__31938\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__7346\ : Odrv4
    port map (
            O => \N__31935\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__7345\ : Odrv4
    port map (
            O => \N__31930\,
            I => \M_this_spr_address_qZ0Z_13\
        );

    \I__7344\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31915\
        );

    \I__7343\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31908\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__31915\,
            I => \N__31905\
        );

    \I__7341\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31902\
        );

    \I__7340\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31899\
        );

    \I__7339\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31895\
        );

    \I__7338\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31892\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31889\
        );

    \I__7336\ : Span4Mux_v
    port map (
            O => \N__31905\,
            I => \N__31884\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__31902\,
            I => \N__31884\
        );

    \I__7334\ : LocalMux
    port map (
            O => \N__31899\,
            I => \N__31881\
        );

    \I__7333\ : InMux
    port map (
            O => \N__31898\,
            I => \N__31878\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__31895\,
            I => \N__31873\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__31892\,
            I => \N__31873\
        );

    \I__7330\ : Span4Mux_h
    port map (
            O => \N__31889\,
            I => \N__31870\
        );

    \I__7329\ : Span4Mux_h
    port map (
            O => \N__31884\,
            I => \N__31867\
        );

    \I__7328\ : Span4Mux_h
    port map (
            O => \N__31881\,
            I => \N__31864\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__31878\,
            I => \N__31861\
        );

    \I__7326\ : Span12Mux_h
    port map (
            O => \N__31873\,
            I => \N__31858\
        );

    \I__7325\ : Span4Mux_h
    port map (
            O => \N__31870\,
            I => \N__31855\
        );

    \I__7324\ : Span4Mux_v
    port map (
            O => \N__31867\,
            I => \N__31850\
        );

    \I__7323\ : Span4Mux_h
    port map (
            O => \N__31864\,
            I => \N__31850\
        );

    \I__7322\ : Span4Mux_h
    port map (
            O => \N__31861\,
            I => \N__31847\
        );

    \I__7321\ : Odrv12
    port map (
            O => \N__31858\,
            I => \M_this_spr_ram_write_en_0_i_1_0\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__31855\,
            I => \M_this_spr_ram_write_en_0_i_1_0\
        );

    \I__7319\ : Odrv4
    port map (
            O => \N__31850\,
            I => \M_this_spr_ram_write_en_0_i_1_0\
        );

    \I__7318\ : Odrv4
    port map (
            O => \N__31847\,
            I => \M_this_spr_ram_write_en_0_i_1_0\
        );

    \I__7317\ : CEMux
    port map (
            O => \N__31838\,
            I => \N__31834\
        );

    \I__7316\ : CEMux
    port map (
            O => \N__31837\,
            I => \N__31831\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31828\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__31831\,
            I => \N__31825\
        );

    \I__7313\ : Span4Mux_v
    port map (
            O => \N__31828\,
            I => \N__31822\
        );

    \I__7312\ : Span4Mux_h
    port map (
            O => \N__31825\,
            I => \N__31819\
        );

    \I__7311\ : Span4Mux_h
    port map (
            O => \N__31822\,
            I => \N__31816\
        );

    \I__7310\ : Span4Mux_h
    port map (
            O => \N__31819\,
            I => \N__31813\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__31816\,
            I => \this_spr_ram.mem_WE_4\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__31813\,
            I => \this_spr_ram.mem_WE_4\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__31808\,
            I => \N__31804\
        );

    \I__7306\ : InMux
    port map (
            O => \N__31807\,
            I => \N__31801\
        );

    \I__7305\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31798\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__31801\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__31798\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\
        );

    \I__7302\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31790\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__31790\,
            I => \this_vga_signals.mult1_un61_sum_axb1_0_1\
        );

    \I__7300\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31784\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__31784\,
            I => \N__31778\
        );

    \I__7298\ : InMux
    port map (
            O => \N__31783\,
            I => \N__31771\
        );

    \I__7297\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31771\
        );

    \I__7296\ : InMux
    port map (
            O => \N__31781\,
            I => \N__31771\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__31778\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__31771\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6\
        );

    \I__7293\ : CascadeMux
    port map (
            O => \N__31766\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_\
        );

    \I__7292\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31760\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__31760\,
            I => \N__31757\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__31757\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_x0\
        );

    \I__7289\ : InMux
    port map (
            O => \N__31754\,
            I => \N__31746\
        );

    \I__7288\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31746\
        );

    \I__7287\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31743\
        );

    \I__7286\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31740\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__31746\,
            I => \N__31732\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__31743\,
            I => \N__31727\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__31740\,
            I => \N__31727\
        );

    \I__7282\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31722\
        );

    \I__7281\ : InMux
    port map (
            O => \N__31738\,
            I => \N__31722\
        );

    \I__7280\ : InMux
    port map (
            O => \N__31737\,
            I => \N__31711\
        );

    \I__7279\ : InMux
    port map (
            O => \N__31736\,
            I => \N__31711\
        );

    \I__7278\ : InMux
    port map (
            O => \N__31735\,
            I => \N__31711\
        );

    \I__7277\ : Span4Mux_h
    port map (
            O => \N__31732\,
            I => \N__31706\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__31727\,
            I => \N__31706\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__31722\,
            I => \N__31703\
        );

    \I__7274\ : InMux
    port map (
            O => \N__31721\,
            I => \N__31700\
        );

    \I__7273\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31693\
        );

    \I__7272\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31693\
        );

    \I__7271\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31693\
        );

    \I__7270\ : LocalMux
    port map (
            O => \N__31711\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns\
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__31706\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns\
        );

    \I__7268\ : Odrv12
    port map (
            O => \N__31703\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__31700\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns\
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__31693\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__31682\,
            I => \this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_\
        );

    \I__7264\ : InMux
    port map (
            O => \N__31679\,
            I => \N__31672\
        );

    \I__7263\ : InMux
    port map (
            O => \N__31678\,
            I => \N__31668\
        );

    \I__7262\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31655\
        );

    \I__7261\ : InMux
    port map (
            O => \N__31676\,
            I => \N__31655\
        );

    \I__7260\ : InMux
    port map (
            O => \N__31675\,
            I => \N__31652\
        );

    \I__7259\ : LocalMux
    port map (
            O => \N__31672\,
            I => \N__31649\
        );

    \I__7258\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31646\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__31668\,
            I => \N__31643\
        );

    \I__7256\ : InMux
    port map (
            O => \N__31667\,
            I => \N__31640\
        );

    \I__7255\ : InMux
    port map (
            O => \N__31666\,
            I => \N__31631\
        );

    \I__7254\ : InMux
    port map (
            O => \N__31665\,
            I => \N__31631\
        );

    \I__7253\ : InMux
    port map (
            O => \N__31664\,
            I => \N__31631\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31663\,
            I => \N__31631\
        );

    \I__7251\ : InMux
    port map (
            O => \N__31662\,
            I => \N__31624\
        );

    \I__7250\ : InMux
    port map (
            O => \N__31661\,
            I => \N__31624\
        );

    \I__7249\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31624\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31619\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__31652\,
            I => \N__31619\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__31649\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__31646\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__31643\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__31640\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__31631\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7241\ : LocalMux
    port map (
            O => \N__31624\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__31619\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1\
        );

    \I__7239\ : InMux
    port map (
            O => \N__31604\,
            I => \N__31601\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__31601\,
            I => \this_vga_signals.g0_2_0_1\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__31598\,
            I => \N__31595\
        );

    \I__7236\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31588\
        );

    \I__7235\ : InMux
    port map (
            O => \N__31594\,
            I => \N__31588\
        );

    \I__7234\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31585\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31588\,
            I => \N__31582\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__31585\,
            I => \this_vga_signals.mult1_un54_sum_axb1_out_0\
        );

    \I__7231\ : Odrv4
    port map (
            O => \N__31582\,
            I => \this_vga_signals.mult1_un54_sum_axb1_out_0\
        );

    \I__7230\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31574\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__31574\,
            I => \N__31569\
        );

    \I__7228\ : InMux
    port map (
            O => \N__31573\,
            I => \N__31566\
        );

    \I__7227\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31563\
        );

    \I__7226\ : Span4Mux_v
    port map (
            O => \N__31569\,
            I => \N__31556\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31556\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31556\
        );

    \I__7223\ : Span4Mux_v
    port map (
            O => \N__31556\,
            I => \N__31553\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__31553\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\
        );

    \I__7221\ : InMux
    port map (
            O => \N__31550\,
            I => \N__31547\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31544\
        );

    \I__7219\ : Sp12to4
    port map (
            O => \N__31544\,
            I => \N__31541\
        );

    \I__7218\ : Span12Mux_h
    port map (
            O => \N__31541\,
            I => \N__31537\
        );

    \I__7217\ : InMux
    port map (
            O => \N__31540\,
            I => \N__31534\
        );

    \I__7216\ : Odrv12
    port map (
            O => \N__31537\,
            I => port_rw_in
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__31534\,
            I => port_rw_in
        );

    \I__7214\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31519\
        );

    \I__7213\ : InMux
    port map (
            O => \N__31528\,
            I => \N__31514\
        );

    \I__7212\ : InMux
    port map (
            O => \N__31527\,
            I => \N__31514\
        );

    \I__7211\ : InMux
    port map (
            O => \N__31526\,
            I => \N__31511\
        );

    \I__7210\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31506\
        );

    \I__7209\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31506\
        );

    \I__7208\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31503\
        );

    \I__7207\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31500\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__31519\,
            I => \N__31489\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__31514\,
            I => \N__31489\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31489\
        );

    \I__7203\ : LocalMux
    port map (
            O => \N__31506\,
            I => \N__31486\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__31503\,
            I => \N__31483\
        );

    \I__7201\ : LocalMux
    port map (
            O => \N__31500\,
            I => \N__31480\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31499\,
            I => \N__31477\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31498\,
            I => \N__31472\
        );

    \I__7198\ : InMux
    port map (
            O => \N__31497\,
            I => \N__31472\
        );

    \I__7197\ : InMux
    port map (
            O => \N__31496\,
            I => \N__31469\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__31489\,
            I => \N__31466\
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__31486\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__31483\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7193\ : Odrv4
    port map (
            O => \N__31480\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__31477\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__31472\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__31469\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7189\ : Odrv4
    port map (
            O => \N__31466\,
            I => \this_vga_signals.mult1_un47_sum_axbxc1\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31448\
        );

    \I__7187\ : LocalMux
    port map (
            O => \N__31448\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9\
        );

    \I__7186\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31442\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__31442\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6\
        );

    \I__7184\ : CascadeMux
    port map (
            O => \N__31439\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_\
        );

    \I__7183\ : CascadeMux
    port map (
            O => \N__31436\,
            I => \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_\
        );

    \I__7182\ : InMux
    port map (
            O => \N__31433\,
            I => \N__31430\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__31430\,
            I => \this_vga_signals.g0_5_5\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__31427\,
            I => \N__31423\
        );

    \I__7179\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31416\
        );

    \I__7178\ : InMux
    port map (
            O => \N__31423\,
            I => \N__31416\
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__31422\,
            I => \N__31413\
        );

    \I__7176\ : CascadeMux
    port map (
            O => \N__31421\,
            I => \N__31402\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__31416\,
            I => \N__31396\
        );

    \I__7174\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31391\
        );

    \I__7173\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31391\
        );

    \I__7172\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31386\
        );

    \I__7171\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31386\
        );

    \I__7170\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31381\
        );

    \I__7169\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31381\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31378\
        );

    \I__7167\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31373\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31373\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31370\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31365\
        );

    \I__7163\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31365\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31399\,
            I => \N__31362\
        );

    \I__7161\ : Span4Mux_v
    port map (
            O => \N__31396\,
            I => \N__31355\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__31391\,
            I => \N__31355\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__31386\,
            I => \N__31355\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__31381\,
            I => \N__31349\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__31378\,
            I => \N__31346\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31339\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__31370\,
            I => \N__31339\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31339\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31336\
        );

    \I__7152\ : Span4Mux_h
    port map (
            O => \N__31355\,
            I => \N__31333\
        );

    \I__7151\ : CascadeMux
    port map (
            O => \N__31354\,
            I => \N__31330\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31353\,
            I => \N__31327\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31324\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__31349\,
            I => \N__31321\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__31346\,
            I => \N__31316\
        );

    \I__7146\ : Span4Mux_v
    port map (
            O => \N__31339\,
            I => \N__31316\
        );

    \I__7145\ : Span4Mux_v
    port map (
            O => \N__31336\,
            I => \N__31311\
        );

    \I__7144\ : Span4Mux_v
    port map (
            O => \N__31333\,
            I => \N__31311\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31330\,
            I => \N__31308\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__31327\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__31324\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__31321\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__31316\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__31311\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7137\ : LocalMux
    port map (
            O => \N__31308\,
            I => \this_vga_signals.M_vcounter_qZ0Z_3\
        );

    \I__7136\ : CascadeMux
    port map (
            O => \N__31295\,
            I => \N__31290\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31294\,
            I => \N__31281\
        );

    \I__7134\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31281\
        );

    \I__7133\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31278\
        );

    \I__7132\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31275\
        );

    \I__7131\ : InMux
    port map (
            O => \N__31288\,
            I => \N__31269\
        );

    \I__7130\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31264\
        );

    \I__7129\ : InMux
    port map (
            O => \N__31286\,
            I => \N__31264\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__31281\,
            I => \N__31261\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__31278\,
            I => \N__31257\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31254\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31274\,
            I => \N__31249\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31273\,
            I => \N__31249\
        );

    \I__7123\ : CascadeMux
    port map (
            O => \N__31272\,
            I => \N__31246\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__31269\,
            I => \N__31243\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31238\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__31261\,
            I => \N__31238\
        );

    \I__7119\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31235\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__31257\,
            I => \N__31230\
        );

    \I__7117\ : Span4Mux_v
    port map (
            O => \N__31254\,
            I => \N__31230\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31227\
        );

    \I__7115\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31223\
        );

    \I__7114\ : Span4Mux_v
    port map (
            O => \N__31243\,
            I => \N__31220\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__31238\,
            I => \N__31217\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__31235\,
            I => \N__31212\
        );

    \I__7111\ : Span4Mux_v
    port map (
            O => \N__31230\,
            I => \N__31212\
        );

    \I__7110\ : Span4Mux_v
    port map (
            O => \N__31227\,
            I => \N__31209\
        );

    \I__7109\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31206\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__31223\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7107\ : Odrv4
    port map (
            O => \N__31220\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7106\ : Odrv4
    port map (
            O => \N__31217\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7105\ : Odrv4
    port map (
            O => \N__31212\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__31209\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__31206\,
            I => \this_vga_signals.M_vcounter_qZ0Z_2\
        );

    \I__7102\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31190\
        );

    \I__7101\ : LocalMux
    port map (
            O => \N__31190\,
            I => \this_vga_signals.N_5_i_1\
        );

    \I__7100\ : InMux
    port map (
            O => \N__31187\,
            I => \N__31184\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__31184\,
            I => \N__31181\
        );

    \I__7098\ : Odrv12
    port map (
            O => \N__31181\,
            I => \this_vga_signals.N_5786_0_0\
        );

    \I__7097\ : InMux
    port map (
            O => \N__31178\,
            I => \N__31175\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__31175\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x0\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__31172\,
            I => \N__31169\
        );

    \I__7094\ : InMux
    port map (
            O => \N__31169\,
            I => \N__31166\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__31166\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_x1\
        );

    \I__7092\ : InMux
    port map (
            O => \N__31163\,
            I => \N__31160\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__31160\,
            I => \N__31156\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31159\,
            I => \N__31153\
        );

    \I__7089\ : Span4Mux_h
    port map (
            O => \N__31156\,
            I => \N__31150\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__31153\,
            I => \this_vga_signals.CO0_0_i_i\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__31150\,
            I => \this_vga_signals.CO0_0_i_i\
        );

    \I__7086\ : InMux
    port map (
            O => \N__31145\,
            I => \N__31142\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31142\,
            I => \N__31139\
        );

    \I__7084\ : Span4Mux_h
    port map (
            O => \N__31139\,
            I => \N__31136\
        );

    \I__7083\ : Odrv4
    port map (
            O => \N__31136\,
            I => \this_vga_signals.N_12_0\
        );

    \I__7082\ : CascadeMux
    port map (
            O => \N__31133\,
            I => \this_vga_signals.N_12_0_cascade_\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31130\,
            I => \N__31126\
        );

    \I__7080\ : InMux
    port map (
            O => \N__31129\,
            I => \N__31123\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__31126\,
            I => \N__31119\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__31123\,
            I => \N__31116\
        );

    \I__7077\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31113\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__31119\,
            I => \N__31110\
        );

    \I__7075\ : Odrv4
    port map (
            O => \N__31116\,
            I => \this_vga_signals.N_7_1_0\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__31113\,
            I => \this_vga_signals.N_7_1_0\
        );

    \I__7073\ : Odrv4
    port map (
            O => \N__31110\,
            I => \this_vga_signals.N_7_1_0\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31103\,
            I => \N__31100\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__31100\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__31097\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31091\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__31091\,
            I => \N__31088\
        );

    \I__7067\ : Span4Mux_h
    port map (
            O => \N__31088\,
            I => \N__31085\
        );

    \I__7066\ : Odrv4
    port map (
            O => \N__31085\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0\
        );

    \I__7065\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31079\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__31079\,
            I => \this_vga_signals.g0_0_1\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31073\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__31073\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_x0\
        );

    \I__7061\ : CascadeMux
    port map (
            O => \N__31070\,
            I => \N__31066\
        );

    \I__7060\ : CascadeMux
    port map (
            O => \N__31069\,
            I => \N__31061\
        );

    \I__7059\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31058\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31053\
        );

    \I__7057\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31053\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31061\,
            I => \N__31050\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__31058\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_1\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__31053\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_1\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__31050\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_1\
        );

    \I__7052\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31040\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__31040\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\
        );

    \I__7050\ : InMux
    port map (
            O => \N__31037\,
            I => \N__31034\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__31034\,
            I => \N__31030\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31033\,
            I => \N__31027\
        );

    \I__7047\ : Span4Mux_h
    port map (
            O => \N__31030\,
            I => \N__31024\
        );

    \I__7046\ : LocalMux
    port map (
            O => \N__31027\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__7045\ : Odrv4
    port map (
            O => \N__31024\,
            I => \this_vga_signals.mult1_un54_sum_axb1\
        );

    \I__7044\ : CascadeMux
    port map (
            O => \N__31019\,
            I => \N__31008\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__31018\,
            I => \N__31005\
        );

    \I__7042\ : CascadeMux
    port map (
            O => \N__31017\,
            I => \N__31002\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__31016\,
            I => \N__30999\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__31015\,
            I => \N__30996\
        );

    \I__7039\ : InMux
    port map (
            O => \N__31014\,
            I => \N__30992\
        );

    \I__7038\ : IoInMux
    port map (
            O => \N__31013\,
            I => \N__30980\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31012\,
            I => \N__30977\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31011\,
            I => \N__30972\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31008\,
            I => \N__30972\
        );

    \I__7034\ : InMux
    port map (
            O => \N__31005\,
            I => \N__30967\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30967\
        );

    \I__7032\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30960\
        );

    \I__7031\ : InMux
    port map (
            O => \N__30996\,
            I => \N__30960\
        );

    \I__7030\ : InMux
    port map (
            O => \N__30995\,
            I => \N__30960\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__30992\,
            I => \N__30957\
        );

    \I__7028\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30954\
        );

    \I__7027\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30951\
        );

    \I__7026\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30946\
        );

    \I__7025\ : InMux
    port map (
            O => \N__30988\,
            I => \N__30946\
        );

    \I__7024\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30939\
        );

    \I__7023\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30939\
        );

    \I__7022\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30939\
        );

    \I__7021\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30936\
        );

    \I__7020\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30933\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__30980\,
            I => \N__30929\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__30977\,
            I => \N__30926\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30915\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__30967\,
            I => \N__30915\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__30960\,
            I => \N__30915\
        );

    \I__7014\ : Span4Mux_h
    port map (
            O => \N__30957\,
            I => \N__30915\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__30954\,
            I => \N__30915\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__30951\,
            I => \N__30912\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__30946\,
            I => \N__30909\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__30939\,
            I => \N__30906\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__30936\,
            I => \N__30901\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30901\
        );

    \I__7007\ : CascadeMux
    port map (
            O => \N__30932\,
            I => \N__30896\
        );

    \I__7006\ : IoSpan4Mux
    port map (
            O => \N__30929\,
            I => \N__30891\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__30926\,
            I => \N__30884\
        );

    \I__7004\ : Span4Mux_h
    port map (
            O => \N__30915\,
            I => \N__30884\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__30912\,
            I => \N__30884\
        );

    \I__7002\ : Span4Mux_v
    port map (
            O => \N__30909\,
            I => \N__30881\
        );

    \I__7001\ : Span4Mux_v
    port map (
            O => \N__30906\,
            I => \N__30878\
        );

    \I__7000\ : Span4Mux_h
    port map (
            O => \N__30901\,
            I => \N__30875\
        );

    \I__6999\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30870\
        );

    \I__6998\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30870\
        );

    \I__6997\ : InMux
    port map (
            O => \N__30896\,
            I => \N__30863\
        );

    \I__6996\ : InMux
    port map (
            O => \N__30895\,
            I => \N__30863\
        );

    \I__6995\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30863\
        );

    \I__6994\ : IoSpan4Mux
    port map (
            O => \N__30891\,
            I => \N__30860\
        );

    \I__6993\ : Span4Mux_v
    port map (
            O => \N__30884\,
            I => \N__30857\
        );

    \I__6992\ : Span4Mux_h
    port map (
            O => \N__30881\,
            I => \N__30852\
        );

    \I__6991\ : Span4Mux_h
    port map (
            O => \N__30878\,
            I => \N__30852\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__30875\,
            I => \N__30849\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__30870\,
            I => \N__30844\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__30863\,
            I => \N__30844\
        );

    \I__6987\ : Sp12to4
    port map (
            O => \N__30860\,
            I => \N__30841\
        );

    \I__6986\ : Span4Mux_h
    port map (
            O => \N__30857\,
            I => \N__30838\
        );

    \I__6985\ : Span4Mux_h
    port map (
            O => \N__30852\,
            I => \N__30835\
        );

    \I__6984\ : Span4Mux_v
    port map (
            O => \N__30849\,
            I => \N__30832\
        );

    \I__6983\ : Span12Mux_v
    port map (
            O => \N__30844\,
            I => \N__30827\
        );

    \I__6982\ : Span12Mux_s9_h
    port map (
            O => \N__30841\,
            I => \N__30827\
        );

    \I__6981\ : Odrv4
    port map (
            O => \N__30838\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6980\ : Odrv4
    port map (
            O => \N__30835\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6979\ : Odrv4
    port map (
            O => \N__30832\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6978\ : Odrv12
    port map (
            O => \N__30827\,
            I => \M_this_reset_cond_out_0\
        );

    \I__6977\ : InMux
    port map (
            O => \N__30818\,
            I => \N__30809\
        );

    \I__6976\ : InMux
    port map (
            O => \N__30817\,
            I => \N__30809\
        );

    \I__6975\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30802\
        );

    \I__6974\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30802\
        );

    \I__6973\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30802\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__30809\,
            I => \N__30795\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__30802\,
            I => \N__30792\
        );

    \I__6970\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30789\
        );

    \I__6969\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30782\
        );

    \I__6968\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30782\
        );

    \I__6967\ : InMux
    port map (
            O => \N__30798\,
            I => \N__30782\
        );

    \I__6966\ : Span4Mux_v
    port map (
            O => \N__30795\,
            I => \N__30778\
        );

    \I__6965\ : Span4Mux_v
    port map (
            O => \N__30792\,
            I => \N__30775\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__30789\,
            I => \N__30772\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30769\
        );

    \I__6962\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30766\
        );

    \I__6961\ : Sp12to4
    port map (
            O => \N__30778\,
            I => \N__30763\
        );

    \I__6960\ : Sp12to4
    port map (
            O => \N__30775\,
            I => \N__30760\
        );

    \I__6959\ : Span4Mux_h
    port map (
            O => \N__30772\,
            I => \N__30757\
        );

    \I__6958\ : Span4Mux_h
    port map (
            O => \N__30769\,
            I => \N__30752\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__30766\,
            I => \N__30752\
        );

    \I__6956\ : Span12Mux_h
    port map (
            O => \N__30763\,
            I => \N__30743\
        );

    \I__6955\ : Span12Mux_h
    port map (
            O => \N__30760\,
            I => \N__30743\
        );

    \I__6954\ : Sp12to4
    port map (
            O => \N__30757\,
            I => \N__30743\
        );

    \I__6953\ : Sp12to4
    port map (
            O => \N__30752\,
            I => \N__30743\
        );

    \I__6952\ : Span12Mux_v
    port map (
            O => \N__30743\,
            I => \N__30740\
        );

    \I__6951\ : Span12Mux_v
    port map (
            O => \N__30740\,
            I => \N__30737\
        );

    \I__6950\ : Odrv12
    port map (
            O => \N__30737\,
            I => rst_n_c
        );

    \I__6949\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30731\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__30731\,
            I => \this_reset_cond.M_stage_qZ0Z_7\
        );

    \I__6947\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30725\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__30725\,
            I => \this_reset_cond.M_stage_qZ0Z_8\
        );

    \I__6945\ : CEMux
    port map (
            O => \N__30722\,
            I => \N__30719\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__30719\,
            I => \N__30715\
        );

    \I__6943\ : CEMux
    port map (
            O => \N__30718\,
            I => \N__30712\
        );

    \I__6942\ : Span4Mux_h
    port map (
            O => \N__30715\,
            I => \N__30709\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__30712\,
            I => \N__30706\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__30709\,
            I => \N__30703\
        );

    \I__6939\ : Span4Mux_h
    port map (
            O => \N__30706\,
            I => \N__30700\
        );

    \I__6938\ : Span4Mux_h
    port map (
            O => \N__30703\,
            I => \N__30697\
        );

    \I__6937\ : Span4Mux_h
    port map (
            O => \N__30700\,
            I => \N__30694\
        );

    \I__6936\ : Odrv4
    port map (
            O => \N__30697\,
            I => \this_spr_ram.mem_WE_10\
        );

    \I__6935\ : Odrv4
    port map (
            O => \N__30694\,
            I => \this_spr_ram.mem_WE_10\
        );

    \I__6934\ : InMux
    port map (
            O => \N__30689\,
            I => \N__30686\
        );

    \I__6933\ : LocalMux
    port map (
            O => \N__30686\,
            I => \this_vga_signals.N_12_0_0\
        );

    \I__6932\ : CascadeMux
    port map (
            O => \N__30683\,
            I => \N__30680\
        );

    \I__6931\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30677\
        );

    \I__6930\ : LocalMux
    port map (
            O => \N__30677\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_4\
        );

    \I__6929\ : InMux
    port map (
            O => \N__30674\,
            I => \N__30671\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__30671\,
            I => \this_vga_signals.M_vcounter_q_fastZ0Z_5\
        );

    \I__6927\ : CascadeMux
    port map (
            O => \N__30668\,
            I => \this_vga_signals.vaddress_c2_cascade_\
        );

    \I__6926\ : InMux
    port map (
            O => \N__30665\,
            I => \N__30662\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30659\
        );

    \I__6924\ : Odrv4
    port map (
            O => \N__30659\,
            I => \this_vga_signals.g1_1\
        );

    \I__6923\ : InMux
    port map (
            O => \N__30656\,
            I => \N__30653\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__30653\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_0\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__30650\,
            I => \this_vga_signals.g0_1_0_cascade_\
        );

    \I__6920\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30644\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30641\
        );

    \I__6918\ : Odrv12
    port map (
            O => \N__30641\,
            I => \this_vga_signals.N_7_1_0_2\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__30638\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__30635\,
            I => \N__30632\
        );

    \I__6915\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30629\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__30629\,
            I => \N__30626\
        );

    \I__6913\ : Odrv4
    port map (
            O => \N__30626\,
            I => \this_vga_signals.g3_1\
        );

    \I__6912\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30620\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__30620\,
            I => \N__30616\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30619\,
            I => \N__30613\
        );

    \I__6909\ : Span4Mux_h
    port map (
            O => \N__30616\,
            I => \N__30610\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__30613\,
            I => \N__30607\
        );

    \I__6907\ : Odrv4
    port map (
            O => \N__30610\,
            I => \this_vga_signals.g1_3\
        );

    \I__6906\ : Odrv12
    port map (
            O => \N__30607\,
            I => \this_vga_signals.g1_3\
        );

    \I__6905\ : InMux
    port map (
            O => \N__30602\,
            I => \N__30599\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__30599\,
            I => \this_vga_signals.N_7_1_0_0\
        );

    \I__6903\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30593\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__30593\,
            I => \this_vga_signals.g0_1_0_0\
        );

    \I__6901\ : InMux
    port map (
            O => \N__30590\,
            I => \N__30587\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__30587\,
            I => \N__30584\
        );

    \I__6899\ : Span4Mux_v
    port map (
            O => \N__30584\,
            I => \N__30577\
        );

    \I__6898\ : InMux
    port map (
            O => \N__30583\,
            I => \N__30572\
        );

    \I__6897\ : InMux
    port map (
            O => \N__30582\,
            I => \N__30572\
        );

    \I__6896\ : InMux
    port map (
            O => \N__30581\,
            I => \N__30569\
        );

    \I__6895\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30566\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__30577\,
            I => \N__30554\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__30572\,
            I => \N__30551\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__30569\,
            I => \N__30548\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__30566\,
            I => \N__30545\
        );

    \I__6890\ : InMux
    port map (
            O => \N__30565\,
            I => \N__30538\
        );

    \I__6889\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30538\
        );

    \I__6888\ : InMux
    port map (
            O => \N__30563\,
            I => \N__30538\
        );

    \I__6887\ : InMux
    port map (
            O => \N__30562\,
            I => \N__30531\
        );

    \I__6886\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30531\
        );

    \I__6885\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30531\
        );

    \I__6884\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30524\
        );

    \I__6883\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30524\
        );

    \I__6882\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30524\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__30554\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6880\ : Odrv4
    port map (
            O => \N__30551\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6879\ : Odrv4
    port map (
            O => \N__30548\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__30545\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__30538\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__30531\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__30524\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns\
        );

    \I__6874\ : InMux
    port map (
            O => \N__30509\,
            I => \N__30506\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__30506\,
            I => \this_vga_signals.g1_0\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__30503\,
            I => \N__30495\
        );

    \I__6871\ : CascadeMux
    port map (
            O => \N__30502\,
            I => \N__30492\
        );

    \I__6870\ : InMux
    port map (
            O => \N__30501\,
            I => \N__30489\
        );

    \I__6869\ : InMux
    port map (
            O => \N__30500\,
            I => \N__30481\
        );

    \I__6868\ : InMux
    port map (
            O => \N__30499\,
            I => \N__30481\
        );

    \I__6867\ : CascadeMux
    port map (
            O => \N__30498\,
            I => \N__30478\
        );

    \I__6866\ : InMux
    port map (
            O => \N__30495\,
            I => \N__30475\
        );

    \I__6865\ : InMux
    port map (
            O => \N__30492\,
            I => \N__30472\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__30489\,
            I => \N__30469\
        );

    \I__6863\ : InMux
    port map (
            O => \N__30488\,
            I => \N__30466\
        );

    \I__6862\ : CascadeMux
    port map (
            O => \N__30487\,
            I => \N__30463\
        );

    \I__6861\ : CascadeMux
    port map (
            O => \N__30486\,
            I => \N__30460\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__30481\,
            I => \N__30457\
        );

    \I__6859\ : InMux
    port map (
            O => \N__30478\,
            I => \N__30454\
        );

    \I__6858\ : LocalMux
    port map (
            O => \N__30475\,
            I => \N__30449\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30449\
        );

    \I__6856\ : Span4Mux_v
    port map (
            O => \N__30469\,
            I => \N__30444\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30444\
        );

    \I__6854\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30439\
        );

    \I__6853\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30439\
        );

    \I__6852\ : Odrv12
    port map (
            O => \N__30457\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__30454\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6850\ : Odrv4
    port map (
            O => \N__30449\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__30444\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__30439\,
            I => \this_vga_signals.mult1_un54_sum_c2_0\
        );

    \I__6847\ : InMux
    port map (
            O => \N__30428\,
            I => \N__30425\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__30425\,
            I => \this_vga_signals.g0_29_1\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__30422\,
            I => \this_vga_signals.g1_0_cascade_\
        );

    \I__6844\ : CascadeMux
    port map (
            O => \N__30419\,
            I => \N__30414\
        );

    \I__6843\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30409\
        );

    \I__6842\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30404\
        );

    \I__6841\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30404\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__30413\,
            I => \N__30400\
        );

    \I__6839\ : CascadeMux
    port map (
            O => \N__30412\,
            I => \N__30394\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__30409\,
            I => \N__30389\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__30404\,
            I => \N__30386\
        );

    \I__6836\ : InMux
    port map (
            O => \N__30403\,
            I => \N__30383\
        );

    \I__6835\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30378\
        );

    \I__6834\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30378\
        );

    \I__6833\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30371\
        );

    \I__6832\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30371\
        );

    \I__6831\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30371\
        );

    \I__6830\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30366\
        );

    \I__6829\ : InMux
    port map (
            O => \N__30392\,
            I => \N__30366\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__30389\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__30386\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__30383\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__30378\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__30371\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__30366\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0
        );

    \I__6822\ : InMux
    port map (
            O => \N__30353\,
            I => \N__30350\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__30350\,
            I => \this_vga_signals.g0_3\
        );

    \I__6820\ : InMux
    port map (
            O => \N__30347\,
            I => \N__30344\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30344\,
            I => \N__30341\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__30341\,
            I => \this_reset_cond.M_stage_qZ0Z_6\
        );

    \I__6817\ : CascadeMux
    port map (
            O => \N__30338\,
            I => \N__30335\
        );

    \I__6816\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30332\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__30332\,
            I => \N__30329\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__30329\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__30326\,
            I => \this_vga_signals.g0_2_0_0_cascade_\
        );

    \I__6812\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30320\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__30320\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_4\
        );

    \I__6810\ : InMux
    port map (
            O => \N__30317\,
            I => \N__30314\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__30314\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0\
        );

    \I__6808\ : CascadeMux
    port map (
            O => \N__30311\,
            I => \N__30308\
        );

    \I__6807\ : InMux
    port map (
            O => \N__30308\,
            I => \N__30305\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__30305\,
            I => \this_vga_signals.g0_6_0\
        );

    \I__6805\ : CascadeMux
    port map (
            O => \N__30302\,
            I => \N__30299\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30296\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__30296\,
            I => \this_vga_signals.g0_0_0_1\
        );

    \I__6802\ : InMux
    port map (
            O => \N__30293\,
            I => \N__30290\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30290\,
            I => \this_vga_signals.g0_5_5_N_2L1\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__30287\,
            I => \N__30284\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30272\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30269\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30282\,
            I => \N__30266\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30281\,
            I => \N__30261\
        );

    \I__6795\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30261\
        );

    \I__6794\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30254\
        );

    \I__6793\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30254\
        );

    \I__6792\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30254\
        );

    \I__6791\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30249\
        );

    \I__6790\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30249\
        );

    \I__6789\ : LocalMux
    port map (
            O => \N__30272\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__30269\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__30266\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__30261\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__30254\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__30249\,
            I => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0
        );

    \I__6783\ : InMux
    port map (
            O => \N__30236\,
            I => \N__30233\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__30233\,
            I => \this_vga_signals.g0_5_0\
        );

    \I__6781\ : CascadeMux
    port map (
            O => \N__30230\,
            I => \N__30224\
        );

    \I__6780\ : InMux
    port map (
            O => \N__30229\,
            I => \N__30214\
        );

    \I__6779\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30214\
        );

    \I__6778\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30211\
        );

    \I__6777\ : InMux
    port map (
            O => \N__30224\,
            I => \N__30204\
        );

    \I__6776\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30204\
        );

    \I__6775\ : InMux
    port map (
            O => \N__30222\,
            I => \N__30204\
        );

    \I__6774\ : InMux
    port map (
            O => \N__30221\,
            I => \N__30197\
        );

    \I__6773\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30197\
        );

    \I__6772\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30197\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__30214\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__6770\ : LocalMux
    port map (
            O => \N__30211\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__30204\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__30197\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3\
        );

    \I__6767\ : CascadeMux
    port map (
            O => \N__30188\,
            I => \this_vga_signals.mult1_un54_sum_c2_0_cascade_\
        );

    \I__6766\ : CascadeMux
    port map (
            O => \N__30185\,
            I => \this_vga_signals.g1_1_0_0_cascade_\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30182\,
            I => \N__30179\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__30179\,
            I => \this_vga_signals.N_20_0\
        );

    \I__6763\ : CascadeMux
    port map (
            O => \N__30176\,
            I => \this_vga_signals.g0_2_0_3_cascade_\
        );

    \I__6762\ : InMux
    port map (
            O => \N__30173\,
            I => \N__30170\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30170\,
            I => \this_vga_signals.g0_0_0_1_0\
        );

    \I__6760\ : InMux
    port map (
            O => \N__30167\,
            I => \N__30164\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__30164\,
            I => \this_vga_signals.g0_0_0\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__30161\,
            I => \this_vga_signals.vaddress_c5_a0_0_cascade_\
        );

    \I__6757\ : CascadeMux
    port map (
            O => \N__30158\,
            I => \this_vga_signals.vaddress_9_cascade_\
        );

    \I__6756\ : CascadeMux
    port map (
            O => \N__30155\,
            I => \this_vga_signals.g1_3_0_cascade_\
        );

    \I__6755\ : CascadeMux
    port map (
            O => \N__30152\,
            I => \this_vga_signals.N_5_0_cascade_\
        );

    \I__6754\ : CascadeMux
    port map (
            O => \N__30149\,
            I => \N__30146\
        );

    \I__6753\ : InMux
    port map (
            O => \N__30146\,
            I => \N__30143\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__30143\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_0_0\
        );

    \I__6751\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30137\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__30137\,
            I => \this_vga_signals.N_4_1\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__30134\,
            I => \this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_\
        );

    \I__6748\ : InMux
    port map (
            O => \N__30131\,
            I => \N__30128\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__30128\,
            I => \this_vga_signals.mult1_un54_sum_c3_x1\
        );

    \I__6746\ : IoInMux
    port map (
            O => \N__30125\,
            I => \N__30122\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30119\
        );

    \I__6744\ : Span4Mux_s2_v
    port map (
            O => \N__30119\,
            I => \N__30116\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__30116\,
            I => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\
        );

    \I__6742\ : CEMux
    port map (
            O => \N__30113\,
            I => \N__30110\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30110\,
            I => \N__30106\
        );

    \I__6740\ : CEMux
    port map (
            O => \N__30109\,
            I => \N__30103\
        );

    \I__6739\ : Span4Mux_v
    port map (
            O => \N__30106\,
            I => \N__30100\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__30103\,
            I => \N__30097\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__30100\,
            I => \N__30092\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__30097\,
            I => \N__30092\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__30092\,
            I => \N__30089\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__30089\,
            I => \this_spr_ram.mem_WE_8\
        );

    \I__6733\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__30083\,
            I => \this_vga_signals.m43_4\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__30080\,
            I => \N__30077\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30074\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__30074\,
            I => \this_vga_signals.vaddress_c3_d_0\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30068\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__30068\,
            I => \N__30065\
        );

    \I__6726\ : Span4Mux_v
    port map (
            O => \N__30065\,
            I => \N__30062\
        );

    \I__6725\ : Odrv4
    port map (
            O => \N__30062\,
            I => \this_vga_signals.g0_1_0_1\
        );

    \I__6724\ : CascadeMux
    port map (
            O => \N__30059\,
            I => \this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_\
        );

    \I__6723\ : CascadeMux
    port map (
            O => \N__30056\,
            I => \this_vga_signals.CO0_0_i_i_cascade_\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__30053\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_\
        );

    \I__6721\ : CascadeMux
    port map (
            O => \N__30050\,
            I => \this_vga_signals.N_5_i_0_cascade_\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30044\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30044\,
            I => \N__30041\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__30041\,
            I => \this_vga_signals.g1_0_0\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__30038\,
            I => \N__30035\
        );

    \I__6716\ : InMux
    port map (
            O => \N__30035\,
            I => \N__30032\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__30032\,
            I => \N__30029\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__30029\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9\
        );

    \I__6713\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30023\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__30023\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2\
        );

    \I__6711\ : CascadeMux
    port map (
            O => \N__30020\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\
        );

    \I__6710\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \N__30014\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30011\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__30011\,
            I => \this_vga_signals.g0_i_x2_1\
        );

    \I__6707\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \this_vga_signals.mult1_un54_sum_c3_x0_cascade_\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__30005\,
            I => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__29999\,
            I => \this_vga_signals.g0_41_N_4L5_1\
        );

    \I__6703\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29993\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__29993\,
            I => \N_6_i\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__29990\,
            I => \this_vga_signals.g0_1_1_cascade_\
        );

    \I__6700\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29984\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__29984\,
            I => \this_vga_signals.mult1_un61_sum_c2_0_0\
        );

    \I__6698\ : InMux
    port map (
            O => \N__29981\,
            I => \N__29978\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__29978\,
            I => \this_vga_signals.g1_4\
        );

    \I__6696\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__29972\,
            I => \this_vga_signals.g1_0_0_0\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \this_vga_signals.g1_0_1_0_cascade_\
        );

    \I__6693\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29963\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__29963\,
            I => \this_vga_signals.N_10\
        );

    \I__6691\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29957\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__29957\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_d_2_0\
        );

    \I__6689\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__6688\ : LocalMux
    port map (
            O => \N__29951\,
            I => \this_vga_signals.g0_0_i_0_1\
        );

    \I__6687\ : CascadeMux
    port map (
            O => \N__29948\,
            I => \this_vga_signals.N_10_i_cascade_\
        );

    \I__6686\ : InMux
    port map (
            O => \N__29945\,
            I => \N__29942\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__29942\,
            I => \N__29939\
        );

    \I__6684\ : Span4Mux_h
    port map (
            O => \N__29939\,
            I => \N__29936\
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__29936\,
            I => \this_vga_signals.g2_1_2\
        );

    \I__6682\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29930\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__29930\,
            I => \this_vga_signals.N_10_i_0\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__29927\,
            I => \this_vga_signals.g0_0_i_0_cascade_\
        );

    \I__6679\ : InMux
    port map (
            O => \N__29924\,
            I => \N__29921\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__29921\,
            I => \this_vga_signals.if_m5_i_0_0\
        );

    \I__6677\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29915\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__29915\,
            I => \this_vga_signals.mult1_un68_sum_c3_0_0_0\
        );

    \I__6675\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29909\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__29909\,
            I => \this_vga_signals.if_N_10_0_0_0\
        );

    \I__6673\ : InMux
    port map (
            O => \N__29906\,
            I => \N__29903\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__29903\,
            I => \this_vga_signals.g0_1_0_3\
        );

    \I__6671\ : InMux
    port map (
            O => \N__29900\,
            I => \N__29897\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__29897\,
            I => \this_vga_signals.g0_1_1_0\
        );

    \I__6669\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\
        );

    \I__6668\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29888\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__29888\,
            I => \this_vga_signals.g0_41_N_3L3_1\
        );

    \I__6666\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29882\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__29882\,
            I => \this_vga_signals.m43_5\
        );

    \I__6664\ : IoInMux
    port map (
            O => \N__29879\,
            I => \N__29876\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__29876\,
            I => \N__29873\
        );

    \I__6662\ : Span4Mux_s3_v
    port map (
            O => \N__29873\,
            I => \N__29870\
        );

    \I__6661\ : Span4Mux_h
    port map (
            O => \N__29870\,
            I => \N__29867\
        );

    \I__6660\ : Span4Mux_v
    port map (
            O => \N__29867\,
            I => \N__29864\
        );

    \I__6659\ : Sp12to4
    port map (
            O => \N__29864\,
            I => \N__29861\
        );

    \I__6658\ : Span12Mux_h
    port map (
            O => \N__29861\,
            I => \N__29858\
        );

    \I__6657\ : Odrv12
    port map (
            O => \N__29858\,
            I => this_vga_signals_vsync_1_i
        );

    \I__6656\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29852\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29849\
        );

    \I__6654\ : Span4Mux_v
    port map (
            O => \N__29849\,
            I => \N__29844\
        );

    \I__6653\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29841\
        );

    \I__6652\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29838\
        );

    \I__6651\ : Span4Mux_h
    port map (
            O => \N__29844\,
            I => \N__29833\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__29841\,
            I => \N__29833\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N_52_0\
        );

    \I__6648\ : Odrv4
    port map (
            O => \N__29833\,
            I => \N_52_0\
        );

    \I__6647\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29825\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__29825\,
            I => \N__29822\
        );

    \I__6645\ : Span4Mux_h
    port map (
            O => \N__29822\,
            I => \N__29818\
        );

    \I__6644\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29815\
        );

    \I__6643\ : Odrv4
    port map (
            O => \N__29818\,
            I => \N_58_0\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__29815\,
            I => \N_58_0\
        );

    \I__6641\ : InMux
    port map (
            O => \N__29810\,
            I => \N__29806\
        );

    \I__6640\ : InMux
    port map (
            O => \N__29809\,
            I => \N__29803\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__29806\,
            I => \N__29798\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29798\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__29798\,
            I => \N__29795\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__29795\,
            I => \this_ppu.line_clk.M_last_qZ0\
        );

    \I__6635\ : CEMux
    port map (
            O => \N__29792\,
            I => \N__29780\
        );

    \I__6634\ : CascadeMux
    port map (
            O => \N__29791\,
            I => \N__29775\
        );

    \I__6633\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29767\
        );

    \I__6632\ : InMux
    port map (
            O => \N__29789\,
            I => \N__29759\
        );

    \I__6631\ : InMux
    port map (
            O => \N__29788\,
            I => \N__29759\
        );

    \I__6630\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29759\
        );

    \I__6629\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29750\
        );

    \I__6628\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29750\
        );

    \I__6627\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29750\
        );

    \I__6626\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29750\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__29780\,
            I => \N__29747\
        );

    \I__6624\ : CascadeMux
    port map (
            O => \N__29779\,
            I => \N__29744\
        );

    \I__6623\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29738\
        );

    \I__6622\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29738\
        );

    \I__6621\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29735\
        );

    \I__6620\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29726\
        );

    \I__6619\ : InMux
    port map (
            O => \N__29772\,
            I => \N__29726\
        );

    \I__6618\ : InMux
    port map (
            O => \N__29771\,
            I => \N__29721\
        );

    \I__6617\ : InMux
    port map (
            O => \N__29770\,
            I => \N__29721\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29718\
        );

    \I__6615\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29715\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__29759\,
            I => \N__29712\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29707\
        );

    \I__6612\ : Span4Mux_h
    port map (
            O => \N__29747\,
            I => \N__29707\
        );

    \I__6611\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29702\
        );

    \I__6610\ : InMux
    port map (
            O => \N__29743\,
            I => \N__29702\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__29738\,
            I => \N__29699\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__29735\,
            I => \N__29696\
        );

    \I__6607\ : InMux
    port map (
            O => \N__29734\,
            I => \N__29687\
        );

    \I__6606\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29687\
        );

    \I__6605\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29687\
        );

    \I__6604\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29687\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__29726\,
            I => \N__29678\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__29721\,
            I => \N__29678\
        );

    \I__6601\ : Span4Mux_v
    port map (
            O => \N__29718\,
            I => \N__29678\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__29715\,
            I => \N__29678\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__29712\,
            I => \N__29673\
        );

    \I__6598\ : Span4Mux_v
    port map (
            O => \N__29707\,
            I => \N__29673\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__29702\,
            I => \N__29664\
        );

    \I__6596\ : Span4Mux_h
    port map (
            O => \N__29699\,
            I => \N__29664\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__29696\,
            I => \N__29664\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__29687\,
            I => \N__29664\
        );

    \I__6593\ : Span4Mux_h
    port map (
            O => \N__29678\,
            I => \N__29661\
        );

    \I__6592\ : Odrv4
    port map (
            O => \N__29673\,
            I => \this_vga_signals.GZ0Z_424\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__29664\,
            I => \this_vga_signals.GZ0Z_424\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__29661\,
            I => \this_vga_signals.GZ0Z_424\
        );

    \I__6589\ : IoInMux
    port map (
            O => \N__29654\,
            I => \N__29651\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__29651\,
            I => \N__29647\
        );

    \I__6587\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29644\
        );

    \I__6586\ : Span12Mux_s8_v
    port map (
            O => \N__29647\,
            I => \N__29641\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__29644\,
            I => \this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9\
        );

    \I__6584\ : Odrv12
    port map (
            O => \N__29641\,
            I => \this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9\
        );

    \I__6583\ : InMux
    port map (
            O => \N__29636\,
            I => \N__29633\
        );

    \I__6582\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29630\
        );

    \I__6581\ : Sp12to4
    port map (
            O => \N__29630\,
            I => \N__29627\
        );

    \I__6580\ : Span12Mux_v
    port map (
            O => \N__29627\,
            I => \N__29624\
        );

    \I__6579\ : Odrv12
    port map (
            O => \N__29624\,
            I => \this_ppu.oam_cache.mem_1\
        );

    \I__6578\ : CascadeMux
    port map (
            O => \N__29621\,
            I => \this_vga_signals.vvisibility_0_cascade_\
        );

    \I__6577\ : CascadeMux
    port map (
            O => \N__29618\,
            I => \N__29614\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29611\
        );

    \I__6575\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29608\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__29611\,
            I => \N__29602\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__29608\,
            I => \N__29602\
        );

    \I__6572\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29599\
        );

    \I__6571\ : Span12Mux_v
    port map (
            O => \N__29602\,
            I => \N__29595\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__29599\,
            I => \N__29592\
        );

    \I__6569\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29589\
        );

    \I__6568\ : Span12Mux_h
    port map (
            O => \N__29595\,
            I => \N__29586\
        );

    \I__6567\ : Span4Mux_h
    port map (
            O => \N__29592\,
            I => \N__29583\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__29589\,
            I => \this_vga_signals.vvisibility\
        );

    \I__6565\ : Odrv12
    port map (
            O => \N__29586\,
            I => \this_vga_signals.vvisibility\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__29583\,
            I => \this_vga_signals.vvisibility\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \N__29566\
        );

    \I__6562\ : CascadeMux
    port map (
            O => \N__29575\,
            I => \N__29563\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__29574\,
            I => \N__29559\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__29573\,
            I => \N__29556\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__29572\,
            I => \N__29552\
        );

    \I__6558\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29547\
        );

    \I__6557\ : CascadeMux
    port map (
            O => \N__29570\,
            I => \N__29543\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__29569\,
            I => \N__29540\
        );

    \I__6555\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29537\
        );

    \I__6554\ : InMux
    port map (
            O => \N__29563\,
            I => \N__29534\
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__29562\,
            I => \N__29531\
        );

    \I__6552\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29528\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29525\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__29555\,
            I => \N__29522\
        );

    \I__6549\ : InMux
    port map (
            O => \N__29552\,
            I => \N__29519\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__29551\,
            I => \N__29516\
        );

    \I__6547\ : CascadeMux
    port map (
            O => \N__29550\,
            I => \N__29511\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29508\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__29546\,
            I => \N__29505\
        );

    \I__6544\ : InMux
    port map (
            O => \N__29543\,
            I => \N__29502\
        );

    \I__6543\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29499\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__29537\,
            I => \N__29494\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__29534\,
            I => \N__29494\
        );

    \I__6540\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29491\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29486\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__29525\,
            I => \N__29486\
        );

    \I__6537\ : InMux
    port map (
            O => \N__29522\,
            I => \N__29483\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__29519\,
            I => \N__29480\
        );

    \I__6535\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29477\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__29515\,
            I => \N__29474\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__29514\,
            I => \N__29471\
        );

    \I__6532\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29468\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29508\,
            I => \N__29465\
        );

    \I__6530\ : InMux
    port map (
            O => \N__29505\,
            I => \N__29462\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29459\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__29499\,
            I => \N__29454\
        );

    \I__6527\ : Span4Mux_v
    port map (
            O => \N__29494\,
            I => \N__29454\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__29491\,
            I => \N__29449\
        );

    \I__6525\ : Span4Mux_v
    port map (
            O => \N__29486\,
            I => \N__29449\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29445\
        );

    \I__6523\ : Span4Mux_v
    port map (
            O => \N__29480\,
            I => \N__29440\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__29477\,
            I => \N__29440\
        );

    \I__6521\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29437\
        );

    \I__6520\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29434\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__29468\,
            I => \N__29427\
        );

    \I__6518\ : Span4Mux_s2_v
    port map (
            O => \N__29465\,
            I => \N__29427\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29427\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__29459\,
            I => \N__29424\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__29454\,
            I => \N__29421\
        );

    \I__6514\ : Sp12to4
    port map (
            O => \N__29449\,
            I => \N__29418\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__29448\,
            I => \N__29415\
        );

    \I__6512\ : Span4Mux_v
    port map (
            O => \N__29445\,
            I => \N__29412\
        );

    \I__6511\ : Span4Mux_v
    port map (
            O => \N__29440\,
            I => \N__29409\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__29437\,
            I => \N__29402\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__29434\,
            I => \N__29402\
        );

    \I__6508\ : Span4Mux_v
    port map (
            O => \N__29427\,
            I => \N__29402\
        );

    \I__6507\ : Span4Mux_h
    port map (
            O => \N__29424\,
            I => \N__29396\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__29421\,
            I => \N__29396\
        );

    \I__6505\ : Span12Mux_h
    port map (
            O => \N__29418\,
            I => \N__29393\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29390\
        );

    \I__6503\ : Sp12to4
    port map (
            O => \N__29412\,
            I => \N__29385\
        );

    \I__6502\ : Sp12to4
    port map (
            O => \N__29409\,
            I => \N__29385\
        );

    \I__6501\ : Sp12to4
    port map (
            O => \N__29402\,
            I => \N__29382\
        );

    \I__6500\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29379\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__29396\,
            I => \N__29376\
        );

    \I__6498\ : Span12Mux_v
    port map (
            O => \N__29393\,
            I => \N__29373\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__29390\,
            I => \N__29366\
        );

    \I__6496\ : Span12Mux_v
    port map (
            O => \N__29385\,
            I => \N__29366\
        );

    \I__6495\ : Span12Mux_s11_v
    port map (
            O => \N__29382\,
            I => \N__29366\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__29379\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__29376\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6492\ : Odrv12
    port map (
            O => \N__29373\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6491\ : Odrv12
    port map (
            O => \N__29366\,
            I => \M_this_spr_address_qZ0Z_7\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29357\,
            I => \un1_M_this_spr_address_q_cry_6\
        );

    \I__6489\ : CascadeMux
    port map (
            O => \N__29354\,
            I => \N__29345\
        );

    \I__6488\ : CascadeMux
    port map (
            O => \N__29353\,
            I => \N__29342\
        );

    \I__6487\ : CascadeMux
    port map (
            O => \N__29352\,
            I => \N__29337\
        );

    \I__6486\ : CascadeMux
    port map (
            O => \N__29351\,
            I => \N__29334\
        );

    \I__6485\ : CascadeMux
    port map (
            O => \N__29350\,
            I => \N__29331\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__29349\,
            I => \N__29328\
        );

    \I__6483\ : CascadeMux
    port map (
            O => \N__29348\,
            I => \N__29325\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29322\
        );

    \I__6481\ : InMux
    port map (
            O => \N__29342\,
            I => \N__29319\
        );

    \I__6480\ : CascadeMux
    port map (
            O => \N__29341\,
            I => \N__29315\
        );

    \I__6479\ : CascadeMux
    port map (
            O => \N__29340\,
            I => \N__29312\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29337\,
            I => \N__29308\
        );

    \I__6477\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29305\
        );

    \I__6476\ : InMux
    port map (
            O => \N__29331\,
            I => \N__29302\
        );

    \I__6475\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29299\
        );

    \I__6474\ : InMux
    port map (
            O => \N__29325\,
            I => \N__29296\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29293\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__29319\,
            I => \N__29290\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__29318\,
            I => \N__29282\
        );

    \I__6470\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29279\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29276\
        );

    \I__6468\ : CascadeMux
    port map (
            O => \N__29311\,
            I => \N__29273\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29268\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__29305\,
            I => \N__29268\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__29302\,
            I => \N__29265\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29260\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__29296\,
            I => \N__29260\
        );

    \I__6462\ : Span4Mux_v
    port map (
            O => \N__29293\,
            I => \N__29255\
        );

    \I__6461\ : Span4Mux_v
    port map (
            O => \N__29290\,
            I => \N__29255\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__29289\,
            I => \N__29252\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__29288\,
            I => \N__29249\
        );

    \I__6458\ : CascadeMux
    port map (
            O => \N__29287\,
            I => \N__29246\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__29286\,
            I => \N__29243\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__29285\,
            I => \N__29240\
        );

    \I__6455\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29237\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__29279\,
            I => \N__29232\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__29276\,
            I => \N__29232\
        );

    \I__6452\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29229\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__29268\,
            I => \N__29224\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__29265\,
            I => \N__29224\
        );

    \I__6449\ : Span4Mux_v
    port map (
            O => \N__29260\,
            I => \N__29221\
        );

    \I__6448\ : Span4Mux_v
    port map (
            O => \N__29255\,
            I => \N__29218\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29215\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29212\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29209\
        );

    \I__6444\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29206\
        );

    \I__6443\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29203\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__29237\,
            I => \N__29196\
        );

    \I__6441\ : Span4Mux_v
    port map (
            O => \N__29232\,
            I => \N__29196\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__29229\,
            I => \N__29196\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__29224\,
            I => \N__29193\
        );

    \I__6438\ : Span4Mux_h
    port map (
            O => \N__29221\,
            I => \N__29187\
        );

    \I__6437\ : Span4Mux_h
    port map (
            O => \N__29218\,
            I => \N__29187\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__29215\,
            I => \N__29180\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__29212\,
            I => \N__29180\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29180\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__29206\,
            I => \N__29173\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29203\,
            I => \N__29173\
        );

    \I__6431\ : Sp12to4
    port map (
            O => \N__29196\,
            I => \N__29173\
        );

    \I__6430\ : Sp12to4
    port map (
            O => \N__29193\,
            I => \N__29170\
        );

    \I__6429\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29167\
        );

    \I__6428\ : Span4Mux_h
    port map (
            O => \N__29187\,
            I => \N__29164\
        );

    \I__6427\ : Span12Mux_v
    port map (
            O => \N__29180\,
            I => \N__29157\
        );

    \I__6426\ : Span12Mux_v
    port map (
            O => \N__29173\,
            I => \N__29157\
        );

    \I__6425\ : Span12Mux_v
    port map (
            O => \N__29170\,
            I => \N__29157\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__29167\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__29164\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__6422\ : Odrv12
    port map (
            O => \N__29157\,
            I => \M_this_spr_address_qZ0Z_8\
        );

    \I__6421\ : InMux
    port map (
            O => \N__29150\,
            I => \bfn_17_13_0_\
        );

    \I__6420\ : CascadeMux
    port map (
            O => \N__29147\,
            I => \N__29144\
        );

    \I__6419\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29139\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__29143\,
            I => \N__29136\
        );

    \I__6417\ : CascadeMux
    port map (
            O => \N__29142\,
            I => \N__29132\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__29139\,
            I => \N__29129\
        );

    \I__6415\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29126\
        );

    \I__6414\ : CascadeMux
    port map (
            O => \N__29135\,
            I => \N__29123\
        );

    \I__6413\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29117\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__29129\,
            I => \N__29112\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__29126\,
            I => \N__29112\
        );

    \I__6410\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29109\
        );

    \I__6409\ : CascadeMux
    port map (
            O => \N__29122\,
            I => \N__29106\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__29121\,
            I => \N__29102\
        );

    \I__6407\ : CascadeMux
    port map (
            O => \N__29120\,
            I => \N__29095\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29088\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__29112\,
            I => \N__29088\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__29109\,
            I => \N__29088\
        );

    \I__6403\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29085\
        );

    \I__6402\ : CascadeMux
    port map (
            O => \N__29105\,
            I => \N__29082\
        );

    \I__6401\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29077\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__29101\,
            I => \N__29074\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__29100\,
            I => \N__29071\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__29099\,
            I => \N__29068\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__29098\,
            I => \N__29065\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29062\
        );

    \I__6395\ : Span4Mux_v
    port map (
            O => \N__29088\,
            I => \N__29057\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29085\,
            I => \N__29057\
        );

    \I__6393\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29054\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__29081\,
            I => \N__29051\
        );

    \I__6391\ : CascadeMux
    port map (
            O => \N__29080\,
            I => \N__29048\
        );

    \I__6390\ : LocalMux
    port map (
            O => \N__29077\,
            I => \N__29044\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29041\
        );

    \I__6388\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29038\
        );

    \I__6387\ : InMux
    port map (
            O => \N__29068\,
            I => \N__29035\
        );

    \I__6386\ : InMux
    port map (
            O => \N__29065\,
            I => \N__29032\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__29062\,
            I => \N__29029\
        );

    \I__6384\ : Span4Mux_h
    port map (
            O => \N__29057\,
            I => \N__29023\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N__29023\
        );

    \I__6382\ : InMux
    port map (
            O => \N__29051\,
            I => \N__29020\
        );

    \I__6381\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29017\
        );

    \I__6380\ : CascadeMux
    port map (
            O => \N__29047\,
            I => \N__29014\
        );

    \I__6379\ : Span4Mux_v
    port map (
            O => \N__29044\,
            I => \N__29011\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__29041\,
            I => \N__29006\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29038\,
            I => \N__29006\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__29035\,
            I => \N__29003\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__29032\,
            I => \N__29000\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__29029\,
            I => \N__28997\
        );

    \I__6373\ : CascadeMux
    port map (
            O => \N__29028\,
            I => \N__28994\
        );

    \I__6372\ : Span4Mux_v
    port map (
            O => \N__29023\,
            I => \N__28987\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__29020\,
            I => \N__28987\
        );

    \I__6370\ : LocalMux
    port map (
            O => \N__29017\,
            I => \N__28987\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29014\,
            I => \N__28984\
        );

    \I__6368\ : Span4Mux_h
    port map (
            O => \N__29011\,
            I => \N__28981\
        );

    \I__6367\ : Span4Mux_v
    port map (
            O => \N__29006\,
            I => \N__28978\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__29003\,
            I => \N__28975\
        );

    \I__6365\ : Span4Mux_h
    port map (
            O => \N__29000\,
            I => \N__28972\
        );

    \I__6364\ : Sp12to4
    port map (
            O => \N__28997\,
            I => \N__28969\
        );

    \I__6363\ : InMux
    port map (
            O => \N__28994\,
            I => \N__28966\
        );

    \I__6362\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28963\
        );

    \I__6361\ : LocalMux
    port map (
            O => \N__28984\,
            I => \N__28960\
        );

    \I__6360\ : Span4Mux_v
    port map (
            O => \N__28981\,
            I => \N__28954\
        );

    \I__6359\ : Span4Mux_h
    port map (
            O => \N__28978\,
            I => \N__28954\
        );

    \I__6358\ : Sp12to4
    port map (
            O => \N__28975\,
            I => \N__28947\
        );

    \I__6357\ : Sp12to4
    port map (
            O => \N__28972\,
            I => \N__28947\
        );

    \I__6356\ : Span12Mux_s7_v
    port map (
            O => \N__28969\,
            I => \N__28947\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__28966\,
            I => \N__28944\
        );

    \I__6354\ : Sp12to4
    port map (
            O => \N__28963\,
            I => \N__28939\
        );

    \I__6353\ : Sp12to4
    port map (
            O => \N__28960\,
            I => \N__28939\
        );

    \I__6352\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28936\
        );

    \I__6351\ : Span4Mux_h
    port map (
            O => \N__28954\,
            I => \N__28933\
        );

    \I__6350\ : Span12Mux_v
    port map (
            O => \N__28947\,
            I => \N__28930\
        );

    \I__6349\ : Span12Mux_h
    port map (
            O => \N__28944\,
            I => \N__28925\
        );

    \I__6348\ : Span12Mux_h
    port map (
            O => \N__28939\,
            I => \N__28925\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__28936\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__6346\ : Odrv4
    port map (
            O => \N__28933\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__6345\ : Odrv12
    port map (
            O => \N__28930\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__6344\ : Odrv12
    port map (
            O => \N__28925\,
            I => \M_this_spr_address_qZ0Z_9\
        );

    \I__6343\ : InMux
    port map (
            O => \N__28916\,
            I => \un1_M_this_spr_address_q_cry_8\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__28913\,
            I => \N__28908\
        );

    \I__6341\ : CascadeMux
    port map (
            O => \N__28912\,
            I => \N__28904\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__28911\,
            I => \N__28895\
        );

    \I__6339\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28891\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__28907\,
            I => \N__28887\
        );

    \I__6337\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28884\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__28903\,
            I => \N__28881\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__28902\,
            I => \N__28878\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__28901\,
            I => \N__28874\
        );

    \I__6333\ : CascadeMux
    port map (
            O => \N__28900\,
            I => \N__28871\
        );

    \I__6332\ : CascadeMux
    port map (
            O => \N__28899\,
            I => \N__28865\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__28898\,
            I => \N__28862\
        );

    \I__6330\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28859\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__28894\,
            I => \N__28856\
        );

    \I__6328\ : LocalMux
    port map (
            O => \N__28891\,
            I => \N__28853\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__28890\,
            I => \N__28850\
        );

    \I__6326\ : InMux
    port map (
            O => \N__28887\,
            I => \N__28847\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28844\
        );

    \I__6324\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28841\
        );

    \I__6323\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28838\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__28877\,
            I => \N__28835\
        );

    \I__6321\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28832\
        );

    \I__6320\ : InMux
    port map (
            O => \N__28871\,
            I => \N__28829\
        );

    \I__6319\ : CascadeMux
    port map (
            O => \N__28870\,
            I => \N__28826\
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__28869\,
            I => \N__28823\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__28868\,
            I => \N__28820\
        );

    \I__6316\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28817\
        );

    \I__6315\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28814\
        );

    \I__6314\ : LocalMux
    port map (
            O => \N__28859\,
            I => \N__28811\
        );

    \I__6313\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28808\
        );

    \I__6312\ : Span4Mux_v
    port map (
            O => \N__28853\,
            I => \N__28805\
        );

    \I__6311\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28802\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__28847\,
            I => \N__28799\
        );

    \I__6309\ : Span4Mux_v
    port map (
            O => \N__28844\,
            I => \N__28792\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__28841\,
            I => \N__28792\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28792\
        );

    \I__6306\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28789\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__28832\,
            I => \N__28784\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__28829\,
            I => \N__28784\
        );

    \I__6303\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28781\
        );

    \I__6302\ : InMux
    port map (
            O => \N__28823\,
            I => \N__28778\
        );

    \I__6301\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28775\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__28817\,
            I => \N__28772\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28767\
        );

    \I__6298\ : Span4Mux_h
    port map (
            O => \N__28811\,
            I => \N__28767\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28764\
        );

    \I__6296\ : Span4Mux_h
    port map (
            O => \N__28805\,
            I => \N__28757\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__28802\,
            I => \N__28757\
        );

    \I__6294\ : Span4Mux_v
    port map (
            O => \N__28799\,
            I => \N__28757\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__28792\,
            I => \N__28752\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28752\
        );

    \I__6291\ : Span4Mux_v
    port map (
            O => \N__28784\,
            I => \N__28745\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28745\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__28778\,
            I => \N__28745\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__28775\,
            I => \N__28742\
        );

    \I__6287\ : Span4Mux_h
    port map (
            O => \N__28772\,
            I => \N__28735\
        );

    \I__6286\ : Span4Mux_v
    port map (
            O => \N__28767\,
            I => \N__28735\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__28764\,
            I => \N__28735\
        );

    \I__6284\ : Span4Mux_v
    port map (
            O => \N__28757\,
            I => \N__28732\
        );

    \I__6283\ : Span4Mux_s2_v
    port map (
            O => \N__28752\,
            I => \N__28729\
        );

    \I__6282\ : Span4Mux_v
    port map (
            O => \N__28745\,
            I => \N__28726\
        );

    \I__6281\ : Span4Mux_s2_v
    port map (
            O => \N__28742\,
            I => \N__28723\
        );

    \I__6280\ : Span4Mux_h
    port map (
            O => \N__28735\,
            I => \N__28719\
        );

    \I__6279\ : Sp12to4
    port map (
            O => \N__28732\,
            I => \N__28716\
        );

    \I__6278\ : Sp12to4
    port map (
            O => \N__28729\,
            I => \N__28713\
        );

    \I__6277\ : Sp12to4
    port map (
            O => \N__28726\,
            I => \N__28708\
        );

    \I__6276\ : Sp12to4
    port map (
            O => \N__28723\,
            I => \N__28708\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28705\
        );

    \I__6274\ : Span4Mux_h
    port map (
            O => \N__28719\,
            I => \N__28702\
        );

    \I__6273\ : Span12Mux_h
    port map (
            O => \N__28716\,
            I => \N__28699\
        );

    \I__6272\ : Span12Mux_h
    port map (
            O => \N__28713\,
            I => \N__28694\
        );

    \I__6271\ : Span12Mux_h
    port map (
            O => \N__28708\,
            I => \N__28694\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28705\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__28702\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__6268\ : Odrv12
    port map (
            O => \N__28699\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__6267\ : Odrv12
    port map (
            O => \N__28694\,
            I => \M_this_spr_address_qZ0Z_10\
        );

    \I__6266\ : InMux
    port map (
            O => \N__28685\,
            I => \un1_M_this_spr_address_q_cry_9\
        );

    \I__6265\ : InMux
    port map (
            O => \N__28682\,
            I => \un1_M_this_spr_address_q_cry_10\
        );

    \I__6264\ : InMux
    port map (
            O => \N__28679\,
            I => \un1_M_this_spr_address_q_cry_11\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28676\,
            I => \un1_M_this_spr_address_q_cry_12\
        );

    \I__6262\ : CascadeMux
    port map (
            O => \N__28673\,
            I => \N__28669\
        );

    \I__6261\ : InMux
    port map (
            O => \N__28672\,
            I => \N__28666\
        );

    \I__6260\ : InMux
    port map (
            O => \N__28669\,
            I => \N__28663\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28658\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__28663\,
            I => \N__28658\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__28658\,
            I => \M_this_spr_ram_write_en_0_i_1\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28651\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28654\,
            I => \N__28648\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28644\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__28648\,
            I => \N__28641\
        );

    \I__6252\ : InMux
    port map (
            O => \N__28647\,
            I => \N__28638\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__28644\,
            I => \N__28635\
        );

    \I__6250\ : Span4Mux_v
    port map (
            O => \N__28641\,
            I => \N__28632\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__28638\,
            I => \N__28629\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__28635\,
            I => \N__28626\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__28632\,
            I => \N__28621\
        );

    \I__6246\ : Span4Mux_h
    port map (
            O => \N__28629\,
            I => \N__28621\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__28626\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__28621\,
            I => \this_vga_signals.M_vcounter_d8\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__28616\,
            I => \N__28607\
        );

    \I__6242\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28604\
        );

    \I__6241\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28597\
        );

    \I__6240\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28597\
        );

    \I__6239\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28597\
        );

    \I__6238\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28593\
        );

    \I__6237\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28590\
        );

    \I__6236\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28587\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28583\
        );

    \I__6234\ : LocalMux
    port map (
            O => \N__28597\,
            I => \N__28580\
        );

    \I__6233\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28577\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28570\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28570\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__28587\,
            I => \N__28570\
        );

    \I__6229\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28564\
        );

    \I__6228\ : Span4Mux_v
    port map (
            O => \N__28583\,
            I => \N__28557\
        );

    \I__6227\ : Span4Mux_h
    port map (
            O => \N__28580\,
            I => \N__28557\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28557\
        );

    \I__6225\ : Span12Mux_h
    port map (
            O => \N__28570\,
            I => \N__28554\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28569\,
            I => \N__28547\
        );

    \I__6223\ : InMux
    port map (
            O => \N__28568\,
            I => \N__28547\
        );

    \I__6222\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28547\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__28564\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__28557\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__6219\ : Odrv12
    port map (
            O => \N__28554\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__28547\,
            I => \this_vga_signals.M_hcounter_d7_0\
        );

    \I__6217\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__28535\,
            I => \N__28531\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__28534\,
            I => \N__28528\
        );

    \I__6214\ : Span4Mux_v
    port map (
            O => \N__28531\,
            I => \N__28525\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28522\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__28525\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__28522\,
            I => \M_this_ctrl_flags_qZ0Z_7\
        );

    \I__6210\ : InMux
    port map (
            O => \N__28517\,
            I => \N__28514\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__28514\,
            I => \N__28511\
        );

    \I__6208\ : Odrv4
    port map (
            O => \N__28511\,
            I => \this_reset_cond.M_stage_qZ0Z_5\
        );

    \I__6207\ : CascadeMux
    port map (
            O => \N__28508\,
            I => \N__28502\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__28507\,
            I => \N__28499\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__28506\,
            I => \N__28496\
        );

    \I__6204\ : CascadeMux
    port map (
            O => \N__28505\,
            I => \N__28492\
        );

    \I__6203\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28487\
        );

    \I__6202\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28484\
        );

    \I__6201\ : InMux
    port map (
            O => \N__28496\,
            I => \N__28481\
        );

    \I__6200\ : CascadeMux
    port map (
            O => \N__28495\,
            I => \N__28478\
        );

    \I__6199\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28474\
        );

    \I__6198\ : CascadeMux
    port map (
            O => \N__28491\,
            I => \N__28471\
        );

    \I__6197\ : CascadeMux
    port map (
            O => \N__28490\,
            I => \N__28466\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__28487\,
            I => \N__28460\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__28484\,
            I => \N__28460\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__28481\,
            I => \N__28456\
        );

    \I__6193\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28453\
        );

    \I__6192\ : CascadeMux
    port map (
            O => \N__28477\,
            I => \N__28450\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28447\
        );

    \I__6190\ : InMux
    port map (
            O => \N__28471\,
            I => \N__28444\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__28470\,
            I => \N__28441\
        );

    \I__6188\ : CascadeMux
    port map (
            O => \N__28469\,
            I => \N__28438\
        );

    \I__6187\ : InMux
    port map (
            O => \N__28466\,
            I => \N__28434\
        );

    \I__6186\ : CascadeMux
    port map (
            O => \N__28465\,
            I => \N__28431\
        );

    \I__6185\ : Span4Mux_v
    port map (
            O => \N__28460\,
            I => \N__28426\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__28459\,
            I => \N__28423\
        );

    \I__6183\ : Span4Mux_s3_v
    port map (
            O => \N__28456\,
            I => \N__28418\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__28453\,
            I => \N__28418\
        );

    \I__6181\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28415\
        );

    \I__6180\ : Span4Mux_s1_v
    port map (
            O => \N__28447\,
            I => \N__28409\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__28444\,
            I => \N__28409\
        );

    \I__6178\ : InMux
    port map (
            O => \N__28441\,
            I => \N__28406\
        );

    \I__6177\ : InMux
    port map (
            O => \N__28438\,
            I => \N__28403\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__28437\,
            I => \N__28400\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28397\
        );

    \I__6174\ : InMux
    port map (
            O => \N__28431\,
            I => \N__28394\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__28430\,
            I => \N__28391\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__28429\,
            I => \N__28388\
        );

    \I__6171\ : Span4Mux_h
    port map (
            O => \N__28426\,
            I => \N__28385\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28382\
        );

    \I__6169\ : Span4Mux_h
    port map (
            O => \N__28418\,
            I => \N__28377\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__28415\,
            I => \N__28377\
        );

    \I__6167\ : CascadeMux
    port map (
            O => \N__28414\,
            I => \N__28374\
        );

    \I__6166\ : Span4Mux_v
    port map (
            O => \N__28409\,
            I => \N__28369\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__28406\,
            I => \N__28369\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__28403\,
            I => \N__28366\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28363\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__28397\,
            I => \N__28358\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__28394\,
            I => \N__28358\
        );

    \I__6160\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28355\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28352\
        );

    \I__6158\ : Span4Mux_h
    port map (
            O => \N__28385\,
            I => \N__28349\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__28382\,
            I => \N__28346\
        );

    \I__6156\ : Span4Mux_v
    port map (
            O => \N__28377\,
            I => \N__28343\
        );

    \I__6155\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28340\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__28369\,
            I => \N__28337\
        );

    \I__6153\ : Span4Mux_v
    port map (
            O => \N__28366\,
            I => \N__28332\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__28363\,
            I => \N__28332\
        );

    \I__6151\ : Span4Mux_v
    port map (
            O => \N__28358\,
            I => \N__28327\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__28355\,
            I => \N__28327\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__28352\,
            I => \N__28324\
        );

    \I__6148\ : Sp12to4
    port map (
            O => \N__28349\,
            I => \N__28319\
        );

    \I__6147\ : Span12Mux_h
    port map (
            O => \N__28346\,
            I => \N__28319\
        );

    \I__6146\ : Sp12to4
    port map (
            O => \N__28343\,
            I => \N__28314\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28314\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__28337\,
            I => \N__28309\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__28332\,
            I => \N__28309\
        );

    \I__6142\ : Span4Mux_h
    port map (
            O => \N__28327\,
            I => \N__28306\
        );

    \I__6141\ : Span4Mux_h
    port map (
            O => \N__28324\,
            I => \N__28303\
        );

    \I__6140\ : Span12Mux_v
    port map (
            O => \N__28319\,
            I => \N__28299\
        );

    \I__6139\ : Span12Mux_h
    port map (
            O => \N__28314\,
            I => \N__28296\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__28309\,
            I => \N__28291\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__28306\,
            I => \N__28291\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__28303\,
            I => \N__28288\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28285\
        );

    \I__6134\ : Odrv12
    port map (
            O => \N__28299\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__6133\ : Odrv12
    port map (
            O => \N__28296\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__6132\ : Odrv4
    port map (
            O => \N__28291\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__6131\ : Odrv4
    port map (
            O => \N__28288\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__28285\,
            I => \M_this_spr_address_qZ0Z_0\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__28274\,
            I => \N__28271\
        );

    \I__6128\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28266\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__28270\,
            I => \N__28263\
        );

    \I__6126\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28258\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28254\
        );

    \I__6124\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28251\
        );

    \I__6123\ : CascadeMux
    port map (
            O => \N__28262\,
            I => \N__28248\
        );

    \I__6122\ : CascadeMux
    port map (
            O => \N__28261\,
            I => \N__28244\
        );

    \I__6121\ : InMux
    port map (
            O => \N__28258\,
            I => \N__28240\
        );

    \I__6120\ : CascadeMux
    port map (
            O => \N__28257\,
            I => \N__28237\
        );

    \I__6119\ : Span4Mux_s3_v
    port map (
            O => \N__28254\,
            I => \N__28230\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28230\
        );

    \I__6117\ : InMux
    port map (
            O => \N__28248\,
            I => \N__28227\
        );

    \I__6116\ : CascadeMux
    port map (
            O => \N__28247\,
            I => \N__28224\
        );

    \I__6115\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28220\
        );

    \I__6114\ : CascadeMux
    port map (
            O => \N__28243\,
            I => \N__28217\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__28240\,
            I => \N__28214\
        );

    \I__6112\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28211\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__28236\,
            I => \N__28208\
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__28235\,
            I => \N__28204\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__28230\,
            I => \N__28198\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__28227\,
            I => \N__28198\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28195\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__28223\,
            I => \N__28192\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__28220\,
            I => \N__28188\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28217\,
            I => \N__28185\
        );

    \I__6103\ : Span4Mux_s3_v
    port map (
            O => \N__28214\,
            I => \N__28179\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__28211\,
            I => \N__28179\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28208\,
            I => \N__28176\
        );

    \I__6100\ : CascadeMux
    port map (
            O => \N__28207\,
            I => \N__28173\
        );

    \I__6099\ : InMux
    port map (
            O => \N__28204\,
            I => \N__28170\
        );

    \I__6098\ : CascadeMux
    port map (
            O => \N__28203\,
            I => \N__28167\
        );

    \I__6097\ : Span4Mux_v
    port map (
            O => \N__28198\,
            I => \N__28162\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28162\
        );

    \I__6095\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28159\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__28191\,
            I => \N__28156\
        );

    \I__6093\ : Span4Mux_v
    port map (
            O => \N__28188\,
            I => \N__28151\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__28185\,
            I => \N__28151\
        );

    \I__6091\ : CascadeMux
    port map (
            O => \N__28184\,
            I => \N__28148\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__28179\,
            I => \N__28143\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28143\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28140\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28137\
        );

    \I__6086\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28134\
        );

    \I__6085\ : Span4Mux_h
    port map (
            O => \N__28162\,
            I => \N__28129\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__28159\,
            I => \N__28129\
        );

    \I__6083\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28126\
        );

    \I__6082\ : Span4Mux_v
    port map (
            O => \N__28151\,
            I => \N__28122\
        );

    \I__6081\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28119\
        );

    \I__6080\ : Span4Mux_v
    port map (
            O => \N__28143\,
            I => \N__28114\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__28140\,
            I => \N__28114\
        );

    \I__6078\ : Span4Mux_v
    port map (
            O => \N__28137\,
            I => \N__28105\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__28134\,
            I => \N__28105\
        );

    \I__6076\ : Span4Mux_v
    port map (
            O => \N__28129\,
            I => \N__28105\
        );

    \I__6075\ : LocalMux
    port map (
            O => \N__28126\,
            I => \N__28105\
        );

    \I__6074\ : CascadeMux
    port map (
            O => \N__28125\,
            I => \N__28102\
        );

    \I__6073\ : Span4Mux_h
    port map (
            O => \N__28122\,
            I => \N__28099\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__28119\,
            I => \N__28096\
        );

    \I__6071\ : Span4Mux_h
    port map (
            O => \N__28114\,
            I => \N__28093\
        );

    \I__6070\ : Span4Mux_v
    port map (
            O => \N__28105\,
            I => \N__28090\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28087\
        );

    \I__6068\ : Sp12to4
    port map (
            O => \N__28099\,
            I => \N__28082\
        );

    \I__6067\ : Span12Mux_s11_h
    port map (
            O => \N__28096\,
            I => \N__28082\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__28093\,
            I => \N__28079\
        );

    \I__6065\ : Sp12to4
    port map (
            O => \N__28090\,
            I => \N__28074\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28087\,
            I => \N__28074\
        );

    \I__6063\ : Span12Mux_v
    port map (
            O => \N__28082\,
            I => \N__28066\
        );

    \I__6062\ : Sp12to4
    port map (
            O => \N__28079\,
            I => \N__28066\
        );

    \I__6061\ : Span12Mux_s8_h
    port map (
            O => \N__28074\,
            I => \N__28066\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28063\
        );

    \I__6059\ : Odrv12
    port map (
            O => \N__28066\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28063\,
            I => \M_this_spr_address_qZ0Z_1\
        );

    \I__6057\ : InMux
    port map (
            O => \N__28058\,
            I => \un1_M_this_spr_address_q_cry_0\
        );

    \I__6056\ : CascadeMux
    port map (
            O => \N__28055\,
            I => \N__28045\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__28054\,
            I => \N__28042\
        );

    \I__6054\ : CascadeMux
    port map (
            O => \N__28053\,
            I => \N__28038\
        );

    \I__6053\ : CascadeMux
    port map (
            O => \N__28052\,
            I => \N__28033\
        );

    \I__6052\ : CascadeMux
    port map (
            O => \N__28051\,
            I => \N__28028\
        );

    \I__6051\ : CascadeMux
    port map (
            O => \N__28050\,
            I => \N__28025\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__28049\,
            I => \N__28022\
        );

    \I__6049\ : CascadeMux
    port map (
            O => \N__28048\,
            I => \N__28019\
        );

    \I__6048\ : InMux
    port map (
            O => \N__28045\,
            I => \N__28016\
        );

    \I__6047\ : InMux
    port map (
            O => \N__28042\,
            I => \N__28013\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__28041\,
            I => \N__28010\
        );

    \I__6045\ : InMux
    port map (
            O => \N__28038\,
            I => \N__28007\
        );

    \I__6044\ : CascadeMux
    port map (
            O => \N__28037\,
            I => \N__28001\
        );

    \I__6043\ : CascadeMux
    port map (
            O => \N__28036\,
            I => \N__27998\
        );

    \I__6042\ : InMux
    port map (
            O => \N__28033\,
            I => \N__27995\
        );

    \I__6041\ : CascadeMux
    port map (
            O => \N__28032\,
            I => \N__27992\
        );

    \I__6040\ : CascadeMux
    port map (
            O => \N__28031\,
            I => \N__27989\
        );

    \I__6039\ : InMux
    port map (
            O => \N__28028\,
            I => \N__27986\
        );

    \I__6038\ : InMux
    port map (
            O => \N__28025\,
            I => \N__27983\
        );

    \I__6037\ : InMux
    port map (
            O => \N__28022\,
            I => \N__27980\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28019\,
            I => \N__27977\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__27974\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__27971\
        );

    \I__6033\ : InMux
    port map (
            O => \N__28010\,
            I => \N__27968\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__28007\,
            I => \N__27965\
        );

    \I__6031\ : CascadeMux
    port map (
            O => \N__28006\,
            I => \N__27962\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__28005\,
            I => \N__27959\
        );

    \I__6029\ : CascadeMux
    port map (
            O => \N__28004\,
            I => \N__27956\
        );

    \I__6028\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27953\
        );

    \I__6027\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27950\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27947\
        );

    \I__6025\ : InMux
    port map (
            O => \N__27992\,
            I => \N__27944\
        );

    \I__6024\ : InMux
    port map (
            O => \N__27989\,
            I => \N__27941\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__27986\,
            I => \N__27938\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__27983\,
            I => \N__27935\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__27980\,
            I => \N__27932\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__27977\,
            I => \N__27929\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__27974\,
            I => \N__27926\
        );

    \I__6018\ : Span4Mux_h
    port map (
            O => \N__27971\,
            I => \N__27923\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__27968\,
            I => \N__27920\
        );

    \I__6016\ : Span4Mux_h
    port map (
            O => \N__27965\,
            I => \N__27917\
        );

    \I__6015\ : InMux
    port map (
            O => \N__27962\,
            I => \N__27914\
        );

    \I__6014\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27911\
        );

    \I__6013\ : InMux
    port map (
            O => \N__27956\,
            I => \N__27908\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__27953\,
            I => \N__27905\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__27950\,
            I => \N__27898\
        );

    \I__6010\ : Span4Mux_v
    port map (
            O => \N__27947\,
            I => \N__27898\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27898\
        );

    \I__6008\ : LocalMux
    port map (
            O => \N__27941\,
            I => \N__27893\
        );

    \I__6007\ : Span4Mux_v
    port map (
            O => \N__27938\,
            I => \N__27893\
        );

    \I__6006\ : Span4Mux_h
    port map (
            O => \N__27935\,
            I => \N__27890\
        );

    \I__6005\ : Span4Mux_h
    port map (
            O => \N__27932\,
            I => \N__27885\
        );

    \I__6004\ : Span4Mux_h
    port map (
            O => \N__27929\,
            I => \N__27885\
        );

    \I__6003\ : Span4Mux_v
    port map (
            O => \N__27926\,
            I => \N__27882\
        );

    \I__6002\ : Span4Mux_v
    port map (
            O => \N__27923\,
            I => \N__27879\
        );

    \I__6001\ : Span4Mux_h
    port map (
            O => \N__27920\,
            I => \N__27874\
        );

    \I__6000\ : Span4Mux_v
    port map (
            O => \N__27917\,
            I => \N__27874\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__27914\,
            I => \N__27871\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__27911\,
            I => \N__27868\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__27908\,
            I => \N__27865\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__27905\,
            I => \N__27860\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__27898\,
            I => \N__27860\
        );

    \I__5994\ : Span4Mux_h
    port map (
            O => \N__27893\,
            I => \N__27854\
        );

    \I__5993\ : Span4Mux_v
    port map (
            O => \N__27890\,
            I => \N__27854\
        );

    \I__5992\ : Sp12to4
    port map (
            O => \N__27885\,
            I => \N__27851\
        );

    \I__5991\ : Sp12to4
    port map (
            O => \N__27882\,
            I => \N__27844\
        );

    \I__5990\ : Sp12to4
    port map (
            O => \N__27879\,
            I => \N__27844\
        );

    \I__5989\ : Sp12to4
    port map (
            O => \N__27874\,
            I => \N__27844\
        );

    \I__5988\ : Span12Mux_h
    port map (
            O => \N__27871\,
            I => \N__27839\
        );

    \I__5987\ : Span12Mux_h
    port map (
            O => \N__27868\,
            I => \N__27839\
        );

    \I__5986\ : Span12Mux_h
    port map (
            O => \N__27865\,
            I => \N__27836\
        );

    \I__5985\ : Span4Mux_h
    port map (
            O => \N__27860\,
            I => \N__27833\
        );

    \I__5984\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27830\
        );

    \I__5983\ : Span4Mux_h
    port map (
            O => \N__27854\,
            I => \N__27827\
        );

    \I__5982\ : Span12Mux_s11_v
    port map (
            O => \N__27851\,
            I => \N__27822\
        );

    \I__5981\ : Span12Mux_v
    port map (
            O => \N__27844\,
            I => \N__27822\
        );

    \I__5980\ : Odrv12
    port map (
            O => \N__27839\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5979\ : Odrv12
    port map (
            O => \N__27836\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5978\ : Odrv4
    port map (
            O => \N__27833\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__27830\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5976\ : Odrv4
    port map (
            O => \N__27827\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5975\ : Odrv12
    port map (
            O => \N__27822\,
            I => \M_this_spr_address_qZ0Z_2\
        );

    \I__5974\ : InMux
    port map (
            O => \N__27809\,
            I => \un1_M_this_spr_address_q_cry_1\
        );

    \I__5973\ : CascadeMux
    port map (
            O => \N__27806\,
            I => \N__27803\
        );

    \I__5972\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27799\
        );

    \I__5971\ : CascadeMux
    port map (
            O => \N__27802\,
            I => \N__27796\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27792\
        );

    \I__5969\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27789\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__27795\,
            I => \N__27786\
        );

    \I__5967\ : Span4Mux_v
    port map (
            O => \N__27792\,
            I => \N__27779\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__27789\,
            I => \N__27779\
        );

    \I__5965\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27776\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__27785\,
            I => \N__27767\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__27784\,
            I => \N__27764\
        );

    \I__5962\ : Span4Mux_h
    port map (
            O => \N__27779\,
            I => \N__27757\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__27776\,
            I => \N__27757\
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__27775\,
            I => \N__27754\
        );

    \I__5959\ : CascadeMux
    port map (
            O => \N__27774\,
            I => \N__27751\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__27773\,
            I => \N__27748\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__27772\,
            I => \N__27745\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__27771\,
            I => \N__27739\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__27770\,
            I => \N__27736\
        );

    \I__5954\ : InMux
    port map (
            O => \N__27767\,
            I => \N__27733\
        );

    \I__5953\ : InMux
    port map (
            O => \N__27764\,
            I => \N__27730\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__27763\,
            I => \N__27727\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__27762\,
            I => \N__27724\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__27757\,
            I => \N__27721\
        );

    \I__5949\ : InMux
    port map (
            O => \N__27754\,
            I => \N__27718\
        );

    \I__5948\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27715\
        );

    \I__5947\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27712\
        );

    \I__5946\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27709\
        );

    \I__5945\ : CascadeMux
    port map (
            O => \N__27744\,
            I => \N__27706\
        );

    \I__5944\ : CascadeMux
    port map (
            O => \N__27743\,
            I => \N__27703\
        );

    \I__5943\ : CascadeMux
    port map (
            O => \N__27742\,
            I => \N__27700\
        );

    \I__5942\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27697\
        );

    \I__5941\ : InMux
    port map (
            O => \N__27736\,
            I => \N__27694\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__27733\,
            I => \N__27689\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__27730\,
            I => \N__27689\
        );

    \I__5938\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27686\
        );

    \I__5937\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27683\
        );

    \I__5936\ : Span4Mux_s1_v
    port map (
            O => \N__27721\,
            I => \N__27678\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__27718\,
            I => \N__27678\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27675\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27672\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__27709\,
            I => \N__27669\
        );

    \I__5931\ : InMux
    port map (
            O => \N__27706\,
            I => \N__27666\
        );

    \I__5930\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27663\
        );

    \I__5929\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27660\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27657\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__27694\,
            I => \N__27652\
        );

    \I__5926\ : Span4Mux_v
    port map (
            O => \N__27689\,
            I => \N__27652\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27647\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__27683\,
            I => \N__27647\
        );

    \I__5923\ : Span4Mux_h
    port map (
            O => \N__27678\,
            I => \N__27644\
        );

    \I__5922\ : Span4Mux_h
    port map (
            O => \N__27675\,
            I => \N__27641\
        );

    \I__5921\ : Span4Mux_h
    port map (
            O => \N__27672\,
            I => \N__27638\
        );

    \I__5920\ : Span4Mux_h
    port map (
            O => \N__27669\,
            I => \N__27635\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__27666\,
            I => \N__27632\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__27663\,
            I => \N__27629\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__27660\,
            I => \N__27626\
        );

    \I__5916\ : Span4Mux_v
    port map (
            O => \N__27657\,
            I => \N__27619\
        );

    \I__5915\ : Span4Mux_v
    port map (
            O => \N__27652\,
            I => \N__27619\
        );

    \I__5914\ : Span4Mux_v
    port map (
            O => \N__27647\,
            I => \N__27619\
        );

    \I__5913\ : Sp12to4
    port map (
            O => \N__27644\,
            I => \N__27616\
        );

    \I__5912\ : Sp12to4
    port map (
            O => \N__27641\,
            I => \N__27609\
        );

    \I__5911\ : Sp12to4
    port map (
            O => \N__27638\,
            I => \N__27609\
        );

    \I__5910\ : Sp12to4
    port map (
            O => \N__27635\,
            I => \N__27609\
        );

    \I__5909\ : Span4Mux_v
    port map (
            O => \N__27632\,
            I => \N__27606\
        );

    \I__5908\ : Span4Mux_v
    port map (
            O => \N__27629\,
            I => \N__27601\
        );

    \I__5907\ : Span4Mux_s2_v
    port map (
            O => \N__27626\,
            I => \N__27601\
        );

    \I__5906\ : Span4Mux_h
    port map (
            O => \N__27619\,
            I => \N__27597\
        );

    \I__5905\ : Span12Mux_v
    port map (
            O => \N__27616\,
            I => \N__27592\
        );

    \I__5904\ : Span12Mux_v
    port map (
            O => \N__27609\,
            I => \N__27592\
        );

    \I__5903\ : Sp12to4
    port map (
            O => \N__27606\,
            I => \N__27587\
        );

    \I__5902\ : Sp12to4
    port map (
            O => \N__27601\,
            I => \N__27587\
        );

    \I__5901\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27584\
        );

    \I__5900\ : Span4Mux_h
    port map (
            O => \N__27597\,
            I => \N__27581\
        );

    \I__5899\ : Span12Mux_h
    port map (
            O => \N__27592\,
            I => \N__27576\
        );

    \I__5898\ : Span12Mux_h
    port map (
            O => \N__27587\,
            I => \N__27576\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__27584\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__27581\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5895\ : Odrv12
    port map (
            O => \N__27576\,
            I => \M_this_spr_address_qZ0Z_3\
        );

    \I__5894\ : InMux
    port map (
            O => \N__27569\,
            I => \un1_M_this_spr_address_q_cry_2\
        );

    \I__5893\ : CascadeMux
    port map (
            O => \N__27566\,
            I => \N__27563\
        );

    \I__5892\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27559\
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__27562\,
            I => \N__27556\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__27559\,
            I => \N__27547\
        );

    \I__5889\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27544\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__27555\,
            I => \N__27541\
        );

    \I__5887\ : CascadeMux
    port map (
            O => \N__27554\,
            I => \N__27537\
        );

    \I__5886\ : CascadeMux
    port map (
            O => \N__27553\,
            I => \N__27534\
        );

    \I__5885\ : CascadeMux
    port map (
            O => \N__27552\,
            I => \N__27529\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__27551\,
            I => \N__27526\
        );

    \I__5883\ : CascadeMux
    port map (
            O => \N__27550\,
            I => \N__27522\
        );

    \I__5882\ : Span4Mux_s3_v
    port map (
            O => \N__27547\,
            I => \N__27516\
        );

    \I__5881\ : LocalMux
    port map (
            O => \N__27544\,
            I => \N__27516\
        );

    \I__5880\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27513\
        );

    \I__5879\ : CascadeMux
    port map (
            O => \N__27540\,
            I => \N__27510\
        );

    \I__5878\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27507\
        );

    \I__5877\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27504\
        );

    \I__5876\ : CascadeMux
    port map (
            O => \N__27533\,
            I => \N__27501\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__27532\,
            I => \N__27498\
        );

    \I__5874\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27493\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27490\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__27525\,
            I => \N__27487\
        );

    \I__5871\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27484\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__27521\,
            I => \N__27481\
        );

    \I__5869\ : Span4Mux_v
    port map (
            O => \N__27516\,
            I => \N__27476\
        );

    \I__5868\ : LocalMux
    port map (
            O => \N__27513\,
            I => \N__27476\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27473\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__27507\,
            I => \N__27470\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27467\
        );

    \I__5864\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27464\
        );

    \I__5863\ : InMux
    port map (
            O => \N__27498\,
            I => \N__27460\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__27497\,
            I => \N__27457\
        );

    \I__5861\ : CascadeMux
    port map (
            O => \N__27496\,
            I => \N__27454\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__27493\,
            I => \N__27451\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27448\
        );

    \I__5858\ : InMux
    port map (
            O => \N__27487\,
            I => \N__27445\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__27484\,
            I => \N__27442\
        );

    \I__5856\ : InMux
    port map (
            O => \N__27481\,
            I => \N__27439\
        );

    \I__5855\ : Span4Mux_h
    port map (
            O => \N__27476\,
            I => \N__27434\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__27473\,
            I => \N__27434\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__27470\,
            I => \N__27427\
        );

    \I__5852\ : Span4Mux_h
    port map (
            O => \N__27467\,
            I => \N__27427\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__27464\,
            I => \N__27427\
        );

    \I__5850\ : CascadeMux
    port map (
            O => \N__27463\,
            I => \N__27424\
        );

    \I__5849\ : LocalMux
    port map (
            O => \N__27460\,
            I => \N__27421\
        );

    \I__5848\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27418\
        );

    \I__5847\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27415\
        );

    \I__5846\ : Span4Mux_v
    port map (
            O => \N__27451\,
            I => \N__27410\
        );

    \I__5845\ : Span4Mux_h
    port map (
            O => \N__27448\,
            I => \N__27410\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27407\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__27442\,
            I => \N__27402\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27402\
        );

    \I__5841\ : Span4Mux_v
    port map (
            O => \N__27434\,
            I => \N__27397\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__27427\,
            I => \N__27397\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27394\
        );

    \I__5838\ : Span12Mux_h
    port map (
            O => \N__27421\,
            I => \N__27391\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__27418\,
            I => \N__27388\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__27415\,
            I => \N__27385\
        );

    \I__5835\ : Sp12to4
    port map (
            O => \N__27410\,
            I => \N__27382\
        );

    \I__5834\ : Sp12to4
    port map (
            O => \N__27407\,
            I => \N__27377\
        );

    \I__5833\ : Sp12to4
    port map (
            O => \N__27402\,
            I => \N__27377\
        );

    \I__5832\ : Sp12to4
    port map (
            O => \N__27397\,
            I => \N__27372\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__27394\,
            I => \N__27372\
        );

    \I__5830\ : Span12Mux_v
    port map (
            O => \N__27391\,
            I => \N__27364\
        );

    \I__5829\ : Span12Mux_h
    port map (
            O => \N__27388\,
            I => \N__27364\
        );

    \I__5828\ : Span12Mux_h
    port map (
            O => \N__27385\,
            I => \N__27364\
        );

    \I__5827\ : Span12Mux_v
    port map (
            O => \N__27382\,
            I => \N__27357\
        );

    \I__5826\ : Span12Mux_s11_v
    port map (
            O => \N__27377\,
            I => \N__27357\
        );

    \I__5825\ : Span12Mux_s11_h
    port map (
            O => \N__27372\,
            I => \N__27357\
        );

    \I__5824\ : InMux
    port map (
            O => \N__27371\,
            I => \N__27354\
        );

    \I__5823\ : Odrv12
    port map (
            O => \N__27364\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__5822\ : Odrv12
    port map (
            O => \N__27357\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__27354\,
            I => \M_this_spr_address_qZ0Z_4\
        );

    \I__5820\ : InMux
    port map (
            O => \N__27347\,
            I => \un1_M_this_spr_address_q_cry_3\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__27344\,
            I => \N__27340\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__27343\,
            I => \N__27337\
        );

    \I__5817\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27330\
        );

    \I__5816\ : InMux
    port map (
            O => \N__27337\,
            I => \N__27327\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__27336\,
            I => \N__27324\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__27335\,
            I => \N__27321\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__27334\,
            I => \N__27313\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__27333\,
            I => \N__27309\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27304\
        );

    \I__5810\ : LocalMux
    port map (
            O => \N__27327\,
            I => \N__27304\
        );

    \I__5809\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27301\
        );

    \I__5808\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27298\
        );

    \I__5807\ : CascadeMux
    port map (
            O => \N__27320\,
            I => \N__27295\
        );

    \I__5806\ : CascadeMux
    port map (
            O => \N__27319\,
            I => \N__27292\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__27318\,
            I => \N__27289\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__27317\,
            I => \N__27286\
        );

    \I__5803\ : CascadeMux
    port map (
            O => \N__27316\,
            I => \N__27283\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27277\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__27312\,
            I => \N__27273\
        );

    \I__5800\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27270\
        );

    \I__5799\ : Span4Mux_v
    port map (
            O => \N__27304\,
            I => \N__27263\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__27301\,
            I => \N__27263\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__27298\,
            I => \N__27263\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27260\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27257\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27289\,
            I => \N__27254\
        );

    \I__5793\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27251\
        );

    \I__5792\ : InMux
    port map (
            O => \N__27283\,
            I => \N__27248\
        );

    \I__5791\ : CascadeMux
    port map (
            O => \N__27282\,
            I => \N__27245\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__27281\,
            I => \N__27242\
        );

    \I__5789\ : CascadeMux
    port map (
            O => \N__27280\,
            I => \N__27239\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__27277\,
            I => \N__27236\
        );

    \I__5787\ : CascadeMux
    port map (
            O => \N__27276\,
            I => \N__27233\
        );

    \I__5786\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27230\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__27270\,
            I => \N__27227\
        );

    \I__5784\ : Span4Mux_v
    port map (
            O => \N__27263\,
            I => \N__27222\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__27260\,
            I => \N__27222\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__27257\,
            I => \N__27217\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__27254\,
            I => \N__27217\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__27251\,
            I => \N__27212\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27212\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27245\,
            I => \N__27209\
        );

    \I__5777\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27206\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27239\,
            I => \N__27203\
        );

    \I__5775\ : Span4Mux_v
    port map (
            O => \N__27236\,
            I => \N__27200\
        );

    \I__5774\ : InMux
    port map (
            O => \N__27233\,
            I => \N__27197\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__27230\,
            I => \N__27194\
        );

    \I__5772\ : Span4Mux_v
    port map (
            O => \N__27227\,
            I => \N__27191\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__27222\,
            I => \N__27188\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__27217\,
            I => \N__27183\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__27212\,
            I => \N__27183\
        );

    \I__5768\ : LocalMux
    port map (
            O => \N__27209\,
            I => \N__27175\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__27206\,
            I => \N__27175\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__27203\,
            I => \N__27175\
        );

    \I__5765\ : Sp12to4
    port map (
            O => \N__27200\,
            I => \N__27166\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__27197\,
            I => \N__27166\
        );

    \I__5763\ : Span12Mux_s8_v
    port map (
            O => \N__27194\,
            I => \N__27166\
        );

    \I__5762\ : Sp12to4
    port map (
            O => \N__27191\,
            I => \N__27166\
        );

    \I__5761\ : Sp12to4
    port map (
            O => \N__27188\,
            I => \N__27163\
        );

    \I__5760\ : Sp12to4
    port map (
            O => \N__27183\,
            I => \N__27160\
        );

    \I__5759\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27157\
        );

    \I__5758\ : Span12Mux_s11_v
    port map (
            O => \N__27175\,
            I => \N__27152\
        );

    \I__5757\ : Span12Mux_v
    port map (
            O => \N__27166\,
            I => \N__27152\
        );

    \I__5756\ : Span12Mux_h
    port map (
            O => \N__27163\,
            I => \N__27147\
        );

    \I__5755\ : Span12Mux_h
    port map (
            O => \N__27160\,
            I => \N__27147\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__27157\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5753\ : Odrv12
    port map (
            O => \N__27152\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5752\ : Odrv12
    port map (
            O => \N__27147\,
            I => \M_this_spr_address_qZ0Z_5\
        );

    \I__5751\ : InMux
    port map (
            O => \N__27140\,
            I => \un1_M_this_spr_address_q_cry_4\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__27137\,
            I => \N__27131\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__27136\,
            I => \N__27127\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27124\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__27134\,
            I => \N__27121\
        );

    \I__5746\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27117\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__27130\,
            I => \N__27114\
        );

    \I__5744\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27110\
        );

    \I__5743\ : InMux
    port map (
            O => \N__27124\,
            I => \N__27107\
        );

    \I__5742\ : InMux
    port map (
            O => \N__27121\,
            I => \N__27102\
        );

    \I__5741\ : CascadeMux
    port map (
            O => \N__27120\,
            I => \N__27099\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27096\
        );

    \I__5739\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27093\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__27113\,
            I => \N__27090\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__27110\,
            I => \N__27087\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__27107\,
            I => \N__27084\
        );

    \I__5735\ : CascadeMux
    port map (
            O => \N__27106\,
            I => \N__27080\
        );

    \I__5734\ : CascadeMux
    port map (
            O => \N__27105\,
            I => \N__27076\
        );

    \I__5733\ : LocalMux
    port map (
            O => \N__27102\,
            I => \N__27070\
        );

    \I__5732\ : InMux
    port map (
            O => \N__27099\,
            I => \N__27067\
        );

    \I__5731\ : Span4Mux_s2_v
    port map (
            O => \N__27096\,
            I => \N__27061\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__27093\,
            I => \N__27061\
        );

    \I__5729\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27058\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__27087\,
            I => \N__27055\
        );

    \I__5727\ : Span4Mux_h
    port map (
            O => \N__27084\,
            I => \N__27052\
        );

    \I__5726\ : CascadeMux
    port map (
            O => \N__27083\,
            I => \N__27049\
        );

    \I__5725\ : InMux
    port map (
            O => \N__27080\,
            I => \N__27046\
        );

    \I__5724\ : CascadeMux
    port map (
            O => \N__27079\,
            I => \N__27043\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27040\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__27075\,
            I => \N__27037\
        );

    \I__5721\ : CascadeMux
    port map (
            O => \N__27074\,
            I => \N__27034\
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__27073\,
            I => \N__27030\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__27070\,
            I => \N__27025\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__27067\,
            I => \N__27025\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__27066\,
            I => \N__27022\
        );

    \I__5716\ : Span4Mux_v
    port map (
            O => \N__27061\,
            I => \N__27017\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27058\,
            I => \N__27017\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__27055\,
            I => \N__27014\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__27052\,
            I => \N__27011\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27049\,
            I => \N__27008\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__27046\,
            I => \N__27005\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27002\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__27040\,
            I => \N__26999\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27037\,
            I => \N__26996\
        );

    \I__5707\ : InMux
    port map (
            O => \N__27034\,
            I => \N__26993\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__27033\,
            I => \N__26990\
        );

    \I__5705\ : InMux
    port map (
            O => \N__27030\,
            I => \N__26987\
        );

    \I__5704\ : Span4Mux_v
    port map (
            O => \N__27025\,
            I => \N__26984\
        );

    \I__5703\ : InMux
    port map (
            O => \N__27022\,
            I => \N__26981\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__27017\,
            I => \N__26978\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__27014\,
            I => \N__26975\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__27011\,
            I => \N__26972\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__27008\,
            I => \N__26969\
        );

    \I__5698\ : Span4Mux_h
    port map (
            O => \N__27005\,
            I => \N__26964\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__27002\,
            I => \N__26964\
        );

    \I__5696\ : Span4Mux_v
    port map (
            O => \N__26999\,
            I => \N__26957\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__26996\,
            I => \N__26957\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26957\
        );

    \I__5693\ : InMux
    port map (
            O => \N__26990\,
            I => \N__26954\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__26987\,
            I => \N__26951\
        );

    \I__5691\ : Sp12to4
    port map (
            O => \N__26984\,
            I => \N__26946\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__26981\,
            I => \N__26946\
        );

    \I__5689\ : Span4Mux_h
    port map (
            O => \N__26978\,
            I => \N__26943\
        );

    \I__5688\ : Sp12to4
    port map (
            O => \N__26975\,
            I => \N__26936\
        );

    \I__5687\ : Sp12to4
    port map (
            O => \N__26972\,
            I => \N__26936\
        );

    \I__5686\ : Span12Mux_h
    port map (
            O => \N__26969\,
            I => \N__26936\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__26964\,
            I => \N__26929\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__26957\,
            I => \N__26929\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26929\
        );

    \I__5682\ : Span12Mux_h
    port map (
            O => \N__26951\,
            I => \N__26923\
        );

    \I__5681\ : Span12Mux_h
    port map (
            O => \N__26946\,
            I => \N__26923\
        );

    \I__5680\ : Span4Mux_h
    port map (
            O => \N__26943\,
            I => \N__26920\
        );

    \I__5679\ : Span12Mux_v
    port map (
            O => \N__26936\,
            I => \N__26915\
        );

    \I__5678\ : Sp12to4
    port map (
            O => \N__26929\,
            I => \N__26915\
        );

    \I__5677\ : InMux
    port map (
            O => \N__26928\,
            I => \N__26912\
        );

    \I__5676\ : Odrv12
    port map (
            O => \N__26923\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__26920\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5674\ : Odrv12
    port map (
            O => \N__26915\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__26912\,
            I => \M_this_spr_address_qZ0Z_6\
        );

    \I__5672\ : InMux
    port map (
            O => \N__26903\,
            I => \un1_M_this_spr_address_q_cry_5\
        );

    \I__5671\ : InMux
    port map (
            O => \N__26900\,
            I => \N__26897\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__26897\,
            I => \M_this_data_count_q_cry_11_THRU_CO\
        );

    \I__5669\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26891\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__26891\,
            I => \M_this_data_count_q_s_13\
        );

    \I__5667\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26885\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__26885\,
            I => \M_this_data_count_q_cry_10_THRU_CO\
        );

    \I__5665\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26877\
        );

    \I__5664\ : InMux
    port map (
            O => \N__26881\,
            I => \N__26874\
        );

    \I__5663\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26871\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26868\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__26874\,
            I => \N__26865\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__26871\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__26868\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__26865\,
            I => \M_this_data_count_qZ0Z_7\
        );

    \I__5657\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26855\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__26855\,
            I => \N__26852\
        );

    \I__5655\ : Odrv4
    port map (
            O => \N__26852\,
            I => \this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11\
        );

    \I__5654\ : CascadeMux
    port map (
            O => \N__26849\,
            I => \this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_\
        );

    \I__5653\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26843\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__26843\,
            I => \this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11\
        );

    \I__5651\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26835\
        );

    \I__5650\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26830\
        );

    \I__5649\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26830\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__26835\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__26830\,
            I => \M_this_data_count_qZ0Z_12\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__26825\,
            I => \N__26822\
        );

    \I__5645\ : InMux
    port map (
            O => \N__26822\,
            I => \N__26817\
        );

    \I__5644\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26812\
        );

    \I__5643\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26812\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__26817\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__26812\,
            I => \M_this_data_count_qZ0Z_11\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__26807\,
            I => \N__26803\
        );

    \I__5639\ : InMux
    port map (
            O => \N__26806\,
            I => \N__26800\
        );

    \I__5638\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26797\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__26800\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__26797\,
            I => \M_this_data_count_qZ0Z_13\
        );

    \I__5635\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26788\
        );

    \I__5634\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26785\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__26788\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__26785\,
            I => \M_this_data_count_qZ0Z_10\
        );

    \I__5631\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26777\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__26777\,
            I => \this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11\
        );

    \I__5629\ : CascadeMux
    port map (
            O => \N__26774\,
            I => \N__26771\
        );

    \I__5628\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__26768\,
            I => \N__26765\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__26765\,
            I => \M_this_data_count_q_cry_5_THRU_CO\
        );

    \I__5625\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26741\
        );

    \I__5624\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26741\
        );

    \I__5623\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26741\
        );

    \I__5622\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26741\
        );

    \I__5621\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26730\
        );

    \I__5620\ : InMux
    port map (
            O => \N__26757\,
            I => \N__26730\
        );

    \I__5619\ : InMux
    port map (
            O => \N__26756\,
            I => \N__26730\
        );

    \I__5618\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26730\
        );

    \I__5617\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26730\
        );

    \I__5616\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26721\
        );

    \I__5615\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26721\
        );

    \I__5614\ : InMux
    port map (
            O => \N__26751\,
            I => \N__26721\
        );

    \I__5613\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26721\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__26741\,
            I => \N_685_i\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__26730\,
            I => \N_685_i\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N_685_i\
        );

    \I__5609\ : CascadeMux
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__5608\ : InMux
    port map (
            O => \N__26711\,
            I => \N__26708\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__26708\,
            I => \N__26705\
        );

    \I__5606\ : Sp12to4
    port map (
            O => \N__26705\,
            I => \N__26700\
        );

    \I__5605\ : InMux
    port map (
            O => \N__26704\,
            I => \N__26695\
        );

    \I__5604\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26695\
        );

    \I__5603\ : Odrv12
    port map (
            O => \N__26700\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__26695\,
            I => \M_this_data_count_qZ0Z_6\
        );

    \I__5601\ : InMux
    port map (
            O => \N__26690\,
            I => \N__26687\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__26687\,
            I => \N__26684\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__26684\,
            I => \N__26680\
        );

    \I__5598\ : InMux
    port map (
            O => \N__26683\,
            I => \N__26677\
        );

    \I__5597\ : Span4Mux_v
    port map (
            O => \N__26680\,
            I => \N__26674\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__26677\,
            I => \M_this_ctrl_flags_qZ0Z_5\
        );

    \I__5595\ : Odrv4
    port map (
            O => \N__26674\,
            I => \M_this_ctrl_flags_qZ0Z_5\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26669\,
            I => \N__26663\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26660\
        );

    \I__5592\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26656\
        );

    \I__5591\ : InMux
    port map (
            O => \N__26666\,
            I => \N__26653\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__26663\,
            I => \N__26648\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__26660\,
            I => \N__26648\
        );

    \I__5588\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26645\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__26656\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__26653\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5585\ : Odrv12
    port map (
            O => \N__26648\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__26645\,
            I => \this_vga_signals.M_vcounter_qZ0Z_1\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__26636\,
            I => \this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_\
        );

    \I__5582\ : InMux
    port map (
            O => \N__26633\,
            I => \N__26630\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__26630\,
            I => \this_vga_signals.g0_i_x2_4\
        );

    \I__5580\ : CascadeMux
    port map (
            O => \N__26627\,
            I => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_\
        );

    \I__5579\ : CascadeMux
    port map (
            O => \N__26624\,
            I => \N__26621\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26618\,
            I => \this_vga_signals.N_17_i\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26612\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__26612\,
            I => \M_this_data_count_q_s_10\
        );

    \I__5574\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26606\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__26606\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_11\
        );

    \I__5572\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26600\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26597\
        );

    \I__5570\ : Span12Mux_h
    port map (
            O => \N__26597\,
            I => \N__26594\
        );

    \I__5569\ : Odrv12
    port map (
            O => \N__26594\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_12\
        );

    \I__5568\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26588\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__26588\,
            I => \this_ppu.M_oam_cache_read_data_i_12\
        );

    \I__5566\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26582\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__26582\,
            I => \N__26579\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__26579\,
            I => \N__26576\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__26576\,
            I => \N__26573\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__26573\,
            I => \N__26570\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__26570\,
            I => \this_ppu.oam_cache.mem_8\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__26567\,
            I => \N__26564\
        );

    \I__5559\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__26561\,
            I => \N__26558\
        );

    \I__5557\ : Span4Mux_v
    port map (
            O => \N__26558\,
            I => \N__26555\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__26555\,
            I => \N__26551\
        );

    \I__5555\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26548\
        );

    \I__5554\ : Odrv4
    port map (
            O => \N__26551\,
            I => \this_ppu.M_oam_cache_read_data_8\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__26548\,
            I => \this_ppu.M_oam_cache_read_data_8\
        );

    \I__5552\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26540\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__26540\,
            I => \N__26537\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__26537\,
            I => \N__26532\
        );

    \I__5549\ : InMux
    port map (
            O => \N__26536\,
            I => \N__26529\
        );

    \I__5548\ : InMux
    port map (
            O => \N__26535\,
            I => \N__26526\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__26532\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__26529\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__26526\,
            I => \this_vga_signals.M_vcounter_qZ0Z_0\
        );

    \I__5544\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \this_vga_signals.N_3_1_cascade_\
        );

    \I__5543\ : InMux
    port map (
            O => \N__26516\,
            I => \N__26513\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__26513\,
            I => \N__26510\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__26510\,
            I => \this_vga_signals.g0_41_N_2L1\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__26507\,
            I => \this_vga_signals.g0_41_N_4L5_cascade_\
        );

    \I__5539\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26501\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__26501\,
            I => \this_vga_signals.g0_41_1\
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__26498\,
            I => \N__26495\
        );

    \I__5536\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26492\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__26492\,
            I => \N__26488\
        );

    \I__5534\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26485\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__26488\,
            I => \N__26482\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__26485\,
            I => \N__26475\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__26482\,
            I => \N__26475\
        );

    \I__5530\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26470\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26470\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__26475\,
            I => \N__26463\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__26470\,
            I => \N__26463\
        );

    \I__5526\ : InMux
    port map (
            O => \N__26469\,
            I => \N__26457\
        );

    \I__5525\ : InMux
    port map (
            O => \N__26468\,
            I => \N__26454\
        );

    \I__5524\ : Span4Mux_h
    port map (
            O => \N__26463\,
            I => \N__26451\
        );

    \I__5523\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26444\
        );

    \I__5522\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26444\
        );

    \I__5521\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26444\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__26457\,
            I => \N__26439\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__26454\,
            I => \N__26439\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__26451\,
            I => \M_this_vga_ramdac_en\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__26444\,
            I => \M_this_vga_ramdac_en\
        );

    \I__5516\ : Odrv4
    port map (
            O => \N__26439\,
            I => \M_this_vga_ramdac_en\
        );

    \I__5515\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__26429\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_0_0_1\
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__5512\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__26420\,
            I => \N__26417\
        );

    \I__5510\ : Span4Mux_h
    port map (
            O => \N__26417\,
            I => \N__26414\
        );

    \I__5509\ : Span4Mux_h
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__26411\,
            I => \M_this_vga_signals_address_7\
        );

    \I__5507\ : InMux
    port map (
            O => \N__26408\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_4\
        );

    \I__5506\ : InMux
    port map (
            O => \N__26405\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_5\
        );

    \I__5505\ : InMux
    port map (
            O => \N__26402\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_6\
        );

    \I__5504\ : InMux
    port map (
            O => \N__26399\,
            I => \bfn_16_16_0_\
        );

    \I__5503\ : InMux
    port map (
            O => \N__26396\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_8\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__26390\,
            I => \this_vga_signals.M_vcounter_d7lto9_i_a2_1\
        );

    \I__5500\ : IoInMux
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__26384\,
            I => \N__26381\
        );

    \I__5498\ : Span4Mux_s3_h
    port map (
            O => \N__26381\,
            I => \N__26378\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__26372\,
            I => \N__26369\
        );

    \I__5494\ : Span4Mux_v
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__5493\ : Odrv4
    port map (
            O => \N__26366\,
            I => port_nmib_1_i
        );

    \I__5492\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__26360\,
            I => \this_ppu.M_oam_cache_read_data_i_11\
        );

    \I__5490\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__26351\,
            I => \N__26348\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__5486\ : Odrv4
    port map (
            O => \N__26345\,
            I => \this_ppu.oam_cache.mem_11\
        );

    \I__5485\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__26339\,
            I => \this_reset_cond.M_stage_qZ0Z_3\
        );

    \I__5483\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__26333\,
            I => \this_reset_cond.M_stage_qZ0Z_4\
        );

    \I__5481\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26327\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__26327\,
            I => \this_reset_cond.M_stage_qZ0Z_0\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26324\,
            I => \N__26321\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__26321\,
            I => \N__26318\
        );

    \I__5477\ : Span4Mux_v
    port map (
            O => \N__26318\,
            I => \N__26315\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__26312\,
            I => \N__26309\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__26303\,
            I => \M_this_map_ram_read_data_0\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__26300\,
            I => \N__26291\
        );

    \I__5470\ : CascadeMux
    port map (
            O => \N__26299\,
            I => \N__26286\
        );

    \I__5469\ : CascadeMux
    port map (
            O => \N__26298\,
            I => \N__26283\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__26297\,
            I => \N__26280\
        );

    \I__5467\ : CascadeMux
    port map (
            O => \N__26296\,
            I => \N__26273\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__26295\,
            I => \N__26270\
        );

    \I__5465\ : CascadeMux
    port map (
            O => \N__26294\,
            I => \N__26267\
        );

    \I__5464\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26264\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__26290\,
            I => \N__26260\
        );

    \I__5462\ : CascadeMux
    port map (
            O => \N__26289\,
            I => \N__26257\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26254\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26283\,
            I => \N__26251\
        );

    \I__5459\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26248\
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__26279\,
            I => \N__26245\
        );

    \I__5457\ : CascadeMux
    port map (
            O => \N__26278\,
            I => \N__26242\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__26277\,
            I => \N__26239\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__26276\,
            I => \N__26236\
        );

    \I__5454\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26233\
        );

    \I__5453\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26230\
        );

    \I__5452\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26227\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__26264\,
            I => \N__26224\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__26263\,
            I => \N__26221\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26260\,
            I => \N__26216\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26213\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26210\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__26251\,
            I => \N__26207\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__26248\,
            I => \N__26204\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26245\,
            I => \N__26201\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26198\
        );

    \I__5442\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26195\
        );

    \I__5441\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26192\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26233\,
            I => \N__26189\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26186\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__26227\,
            I => \N__26183\
        );

    \I__5437\ : Span4Mux_v
    port map (
            O => \N__26224\,
            I => \N__26180\
        );

    \I__5436\ : InMux
    port map (
            O => \N__26221\,
            I => \N__26177\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__26220\,
            I => \N__26174\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__26219\,
            I => \N__26171\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26168\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26165\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__26210\,
            I => \N__26162\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__26207\,
            I => \N__26159\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__26204\,
            I => \N__26156\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__26201\,
            I => \N__26153\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26148\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__26195\,
            I => \N__26148\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__26192\,
            I => \N__26141\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__26189\,
            I => \N__26141\
        );

    \I__5423\ : Span4Mux_v
    port map (
            O => \N__26186\,
            I => \N__26141\
        );

    \I__5422\ : Sp12to4
    port map (
            O => \N__26183\,
            I => \N__26138\
        );

    \I__5421\ : Sp12to4
    port map (
            O => \N__26180\,
            I => \N__26133\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__26177\,
            I => \N__26133\
        );

    \I__5419\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26130\
        );

    \I__5418\ : InMux
    port map (
            O => \N__26171\,
            I => \N__26127\
        );

    \I__5417\ : Span4Mux_h
    port map (
            O => \N__26168\,
            I => \N__26124\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__26165\,
            I => \N__26121\
        );

    \I__5415\ : Span4Mux_h
    port map (
            O => \N__26162\,
            I => \N__26118\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__26159\,
            I => \N__26113\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__26156\,
            I => \N__26113\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__26153\,
            I => \N__26106\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__26148\,
            I => \N__26106\
        );

    \I__5410\ : Span4Mux_v
    port map (
            O => \N__26141\,
            I => \N__26106\
        );

    \I__5409\ : Span12Mux_h
    port map (
            O => \N__26138\,
            I => \N__26101\
        );

    \I__5408\ : Span12Mux_h
    port map (
            O => \N__26133\,
            I => \N__26101\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26130\,
            I => \N__26098\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26095\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__26124\,
            I => \N__26090\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__26121\,
            I => \N__26090\
        );

    \I__5403\ : Sp12to4
    port map (
            O => \N__26118\,
            I => \N__26085\
        );

    \I__5402\ : Sp12to4
    port map (
            O => \N__26113\,
            I => \N__26085\
        );

    \I__5401\ : Sp12to4
    port map (
            O => \N__26106\,
            I => \N__26080\
        );

    \I__5400\ : Span12Mux_v
    port map (
            O => \N__26101\,
            I => \N__26080\
        );

    \I__5399\ : Span12Mux_h
    port map (
            O => \N__26098\,
            I => \N__26071\
        );

    \I__5398\ : Span12Mux_h
    port map (
            O => \N__26095\,
            I => \N__26071\
        );

    \I__5397\ : Sp12to4
    port map (
            O => \N__26090\,
            I => \N__26071\
        );

    \I__5396\ : Span12Mux_v
    port map (
            O => \N__26085\,
            I => \N__26071\
        );

    \I__5395\ : Odrv12
    port map (
            O => \N__26080\,
            I => \M_this_ppu_spr_addr_6\
        );

    \I__5394\ : Odrv12
    port map (
            O => \N__26071\,
            I => \M_this_ppu_spr_addr_6\
        );

    \I__5393\ : InMux
    port map (
            O => \N__26066\,
            I => \N__26063\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__5391\ : Sp12to4
    port map (
            O => \N__26060\,
            I => \N__26057\
        );

    \I__5390\ : Span12Mux_v
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__5389\ : Odrv12
    port map (
            O => \N__26054\,
            I => \this_ppu.oam_cache.mem_0\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__26048\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\
        );

    \I__5386\ : InMux
    port map (
            O => \N__26045\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_0\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26042\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_1\
        );

    \I__5384\ : InMux
    port map (
            O => \N__26039\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_2\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26036\,
            I => \this_vga_signals.un1_M_vcounter_q_cry_3\
        );

    \I__5382\ : InMux
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__5380\ : Span4Mux_h
    port map (
            O => \N__26027\,
            I => \N__26024\
        );

    \I__5379\ : Odrv4
    port map (
            O => \N__26024\,
            I => \M_this_data_count_q_cry_3_THRU_CO\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__5377\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26015\,
            I => \N__26010\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26014\,
            I => \N__26005\
        );

    \I__5374\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26005\
        );

    \I__5373\ : Odrv4
    port map (
            O => \N__26010\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__26005\,
            I => \M_this_data_count_qZ0Z_4\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__26000\,
            I => \N__25997\
        );

    \I__5370\ : InMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__5368\ : Odrv12
    port map (
            O => \N__25991\,
            I => \M_this_data_count_q_cry_4_THRU_CO\
        );

    \I__5367\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__25985\,
            I => \N__25980\
        );

    \I__5365\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25975\
        );

    \I__5364\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25975\
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__25980\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__25975\,
            I => \M_this_data_count_qZ0Z_5\
        );

    \I__5361\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25967\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__25967\,
            I => \M_this_data_count_q_cry_8_THRU_CO\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__25964\,
            I => \N__25960\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__25963\,
            I => \N__25956\
        );

    \I__5357\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25953\
        );

    \I__5356\ : InMux
    port map (
            O => \N__25959\,
            I => \N__25948\
        );

    \I__5355\ : InMux
    port map (
            O => \N__25956\,
            I => \N__25948\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__25953\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__25948\,
            I => \M_this_data_count_qZ0Z_9\
        );

    \I__5352\ : InMux
    port map (
            O => \N__25943\,
            I => \N__25938\
        );

    \I__5351\ : InMux
    port map (
            O => \N__25942\,
            I => \N__25933\
        );

    \I__5350\ : InMux
    port map (
            O => \N__25941\,
            I => \N__25930\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__25938\,
            I => \N__25927\
        );

    \I__5348\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25924\
        );

    \I__5347\ : InMux
    port map (
            O => \N__25936\,
            I => \N__25921\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__25933\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__25930\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__5344\ : Odrv4
    port map (
            O => \N__25927\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__25924\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__25921\,
            I => \this_start_data_delay.M_last_qZ0\
        );

    \I__5341\ : CascadeMux
    port map (
            O => \N__25910\,
            I => \N_685_i_cascade_\
        );

    \I__5340\ : CascadeMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__5339\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25900\
        );

    \I__5338\ : InMux
    port map (
            O => \N__25903\,
            I => \N__25896\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__25900\,
            I => \N__25893\
        );

    \I__5336\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25890\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__25896\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__25893\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__25890\,
            I => \M_this_data_count_qZ0Z_2\
        );

    \I__5332\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25879\
        );

    \I__5331\ : InMux
    port map (
            O => \N__25882\,
            I => \N__25875\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__25879\,
            I => \N__25872\
        );

    \I__5329\ : InMux
    port map (
            O => \N__25878\,
            I => \N__25869\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__25875\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__25872\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__25869\,
            I => \M_this_data_count_qZ0Z_1\
        );

    \I__5325\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25857\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__25861\,
            I => \N__25854\
        );

    \I__5323\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25851\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__25857\,
            I => \N__25848\
        );

    \I__5321\ : InMux
    port map (
            O => \N__25854\,
            I => \N__25845\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__25851\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__5319\ : Odrv4
    port map (
            O => \N__25848\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__25845\,
            I => \M_this_data_count_qZ0Z_3\
        );

    \I__5317\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25835\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__25835\,
            I => \N__25830\
        );

    \I__5315\ : InMux
    port map (
            O => \N__25834\,
            I => \N__25825\
        );

    \I__5314\ : InMux
    port map (
            O => \N__25833\,
            I => \N__25825\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__25830\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__25825\,
            I => \M_this_data_count_qZ0Z_0\
        );

    \I__5311\ : InMux
    port map (
            O => \N__25820\,
            I => \N__25817\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__25817\,
            I => \this_reset_cond.M_stage_qZ0Z_1\
        );

    \I__5309\ : InMux
    port map (
            O => \N__25814\,
            I => \M_this_data_count_q_cry_8\
        );

    \I__5308\ : InMux
    port map (
            O => \N__25811\,
            I => \M_this_data_count_q_cry_9\
        );

    \I__5307\ : InMux
    port map (
            O => \N__25808\,
            I => \M_this_data_count_q_cry_10\
        );

    \I__5306\ : IoInMux
    port map (
            O => \N__25805\,
            I => \N__25802\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25792\
        );

    \I__5304\ : SRMux
    port map (
            O => \N__25801\,
            I => \N__25789\
        );

    \I__5303\ : SRMux
    port map (
            O => \N__25800\,
            I => \N__25784\
        );

    \I__5302\ : SRMux
    port map (
            O => \N__25799\,
            I => \N__25781\
        );

    \I__5301\ : SRMux
    port map (
            O => \N__25798\,
            I => \N__25778\
        );

    \I__5300\ : SRMux
    port map (
            O => \N__25797\,
            I => \N__25773\
        );

    \I__5299\ : SRMux
    port map (
            O => \N__25796\,
            I => \N__25770\
        );

    \I__5298\ : SRMux
    port map (
            O => \N__25795\,
            I => \N__25767\
        );

    \I__5297\ : IoSpan4Mux
    port map (
            O => \N__25792\,
            I => \N__25761\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25758\
        );

    \I__5295\ : SRMux
    port map (
            O => \N__25788\,
            I => \N__25755\
        );

    \I__5294\ : SRMux
    port map (
            O => \N__25787\,
            I => \N__25752\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__25784\,
            I => \N__25749\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__25781\,
            I => \N__25744\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__25778\,
            I => \N__25744\
        );

    \I__5290\ : SRMux
    port map (
            O => \N__25777\,
            I => \N__25741\
        );

    \I__5289\ : SRMux
    port map (
            O => \N__25776\,
            I => \N__25738\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25733\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__25770\,
            I => \N__25728\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__25767\,
            I => \N__25728\
        );

    \I__5285\ : SRMux
    port map (
            O => \N__25766\,
            I => \N__25725\
        );

    \I__5284\ : SRMux
    port map (
            O => \N__25765\,
            I => \N__25714\
        );

    \I__5283\ : SRMux
    port map (
            O => \N__25764\,
            I => \N__25711\
        );

    \I__5282\ : Span4Mux_s3_h
    port map (
            O => \N__25761\,
            I => \N__25708\
        );

    \I__5281\ : Span4Mux_s3_v
    port map (
            O => \N__25758\,
            I => \N__25701\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__25755\,
            I => \N__25701\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25701\
        );

    \I__5278\ : Span4Mux_s3_v
    port map (
            O => \N__25749\,
            I => \N__25692\
        );

    \I__5277\ : Span4Mux_s3_v
    port map (
            O => \N__25744\,
            I => \N__25692\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__25741\,
            I => \N__25692\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__25738\,
            I => \N__25692\
        );

    \I__5274\ : SRMux
    port map (
            O => \N__25737\,
            I => \N__25689\
        );

    \I__5273\ : SRMux
    port map (
            O => \N__25736\,
            I => \N__25686\
        );

    \I__5272\ : Span4Mux_s3_v
    port map (
            O => \N__25733\,
            I => \N__25671\
        );

    \I__5271\ : Span4Mux_s3_v
    port map (
            O => \N__25728\,
            I => \N__25671\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__25725\,
            I => \N__25671\
        );

    \I__5269\ : SRMux
    port map (
            O => \N__25724\,
            I => \N__25668\
        );

    \I__5268\ : SRMux
    port map (
            O => \N__25723\,
            I => \N__25665\
        );

    \I__5267\ : SRMux
    port map (
            O => \N__25722\,
            I => \N__25662\
        );

    \I__5266\ : SRMux
    port map (
            O => \N__25721\,
            I => \N__25657\
        );

    \I__5265\ : SRMux
    port map (
            O => \N__25720\,
            I => \N__25654\
        );

    \I__5264\ : SRMux
    port map (
            O => \N__25719\,
            I => \N__25651\
        );

    \I__5263\ : SRMux
    port map (
            O => \N__25718\,
            I => \N__25648\
        );

    \I__5262\ : SRMux
    port map (
            O => \N__25717\,
            I => \N__25645\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__25714\,
            I => \N__25640\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__25711\,
            I => \N__25640\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__25708\,
            I => \N__25629\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__25701\,
            I => \N__25629\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__25692\,
            I => \N__25629\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25689\,
            I => \N__25629\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__25686\,
            I => \N__25629\
        );

    \I__5254\ : SRMux
    port map (
            O => \N__25685\,
            I => \N__25626\
        );

    \I__5253\ : SRMux
    port map (
            O => \N__25684\,
            I => \N__25622\
        );

    \I__5252\ : SRMux
    port map (
            O => \N__25683\,
            I => \N__25619\
        );

    \I__5251\ : IoInMux
    port map (
            O => \N__25682\,
            I => \N__25615\
        );

    \I__5250\ : SRMux
    port map (
            O => \N__25681\,
            I => \N__25612\
        );

    \I__5249\ : SRMux
    port map (
            O => \N__25680\,
            I => \N__25609\
        );

    \I__5248\ : SRMux
    port map (
            O => \N__25679\,
            I => \N__25606\
        );

    \I__5247\ : SRMux
    port map (
            O => \N__25678\,
            I => \N__25603\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__25671\,
            I => \N__25594\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__25668\,
            I => \N__25594\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__25665\,
            I => \N__25589\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__25662\,
            I => \N__25589\
        );

    \I__5242\ : SRMux
    port map (
            O => \N__25661\,
            I => \N__25586\
        );

    \I__5241\ : SRMux
    port map (
            O => \N__25660\,
            I => \N__25583\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25575\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__25654\,
            I => \N__25575\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__25651\,
            I => \N__25570\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25570\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__25645\,
            I => \N__25567\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__25640\,
            I => \N__25560\
        );

    \I__5234\ : Span4Mux_v
    port map (
            O => \N__25629\,
            I => \N__25560\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__25626\,
            I => \N__25560\
        );

    \I__5232\ : SRMux
    port map (
            O => \N__25625\,
            I => \N__25557\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25554\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__25619\,
            I => \N__25551\
        );

    \I__5229\ : SRMux
    port map (
            O => \N__25618\,
            I => \N__25548\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__25615\,
            I => \N__25545\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__25612\,
            I => \N__25538\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__25609\,
            I => \N__25538\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__25606\,
            I => \N__25533\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__25603\,
            I => \N__25533\
        );

    \I__5223\ : SRMux
    port map (
            O => \N__25602\,
            I => \N__25530\
        );

    \I__5222\ : SRMux
    port map (
            O => \N__25601\,
            I => \N__25527\
        );

    \I__5221\ : SRMux
    port map (
            O => \N__25600\,
            I => \N__25524\
        );

    \I__5220\ : SRMux
    port map (
            O => \N__25599\,
            I => \N__25521\
        );

    \I__5219\ : Span4Mux_h
    port map (
            O => \N__25594\,
            I => \N__25516\
        );

    \I__5218\ : Span4Mux_v
    port map (
            O => \N__25589\,
            I => \N__25516\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__25586\,
            I => \N__25510\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__25583\,
            I => \N__25510\
        );

    \I__5215\ : SRMux
    port map (
            O => \N__25582\,
            I => \N__25507\
        );

    \I__5214\ : SRMux
    port map (
            O => \N__25581\,
            I => \N__25504\
        );

    \I__5213\ : SRMux
    port map (
            O => \N__25580\,
            I => \N__25500\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__25575\,
            I => \N__25497\
        );

    \I__5211\ : Span4Mux_v
    port map (
            O => \N__25570\,
            I => \N__25494\
        );

    \I__5210\ : Span4Mux_h
    port map (
            O => \N__25567\,
            I => \N__25487\
        );

    \I__5209\ : Span4Mux_v
    port map (
            O => \N__25560\,
            I => \N__25487\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__25557\,
            I => \N__25487\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__25554\,
            I => \N__25480\
        );

    \I__5206\ : Span4Mux_v
    port map (
            O => \N__25551\,
            I => \N__25480\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__25548\,
            I => \N__25480\
        );

    \I__5204\ : IoSpan4Mux
    port map (
            O => \N__25545\,
            I => \N__25477\
        );

    \I__5203\ : SRMux
    port map (
            O => \N__25544\,
            I => \N__25474\
        );

    \I__5202\ : SRMux
    port map (
            O => \N__25543\,
            I => \N__25471\
        );

    \I__5201\ : Span4Mux_v
    port map (
            O => \N__25538\,
            I => \N__25462\
        );

    \I__5200\ : Span4Mux_v
    port map (
            O => \N__25533\,
            I => \N__25462\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__25530\,
            I => \N__25462\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__25527\,
            I => \N__25462\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25457\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__25521\,
            I => \N__25457\
        );

    \I__5195\ : Span4Mux_v
    port map (
            O => \N__25516\,
            I => \N__25454\
        );

    \I__5194\ : SRMux
    port map (
            O => \N__25515\,
            I => \N__25451\
        );

    \I__5193\ : Span4Mux_v
    port map (
            O => \N__25510\,
            I => \N__25444\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__25507\,
            I => \N__25444\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25444\
        );

    \I__5190\ : SRMux
    port map (
            O => \N__25503\,
            I => \N__25441\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__25500\,
            I => \N__25438\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__25497\,
            I => \N__25431\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__25494\,
            I => \N__25431\
        );

    \I__5186\ : Span4Mux_v
    port map (
            O => \N__25487\,
            I => \N__25431\
        );

    \I__5185\ : Span4Mux_v
    port map (
            O => \N__25480\,
            I => \N__25428\
        );

    \I__5184\ : Span4Mux_s3_h
    port map (
            O => \N__25477\,
            I => \N__25425\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__25474\,
            I => \N__25420\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__25471\,
            I => \N__25420\
        );

    \I__5181\ : Span4Mux_v
    port map (
            O => \N__25462\,
            I => \N__25415\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__25457\,
            I => \N__25415\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__25454\,
            I => \N__25406\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__25451\,
            I => \N__25406\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__25444\,
            I => \N__25406\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25406\
        );

    \I__5175\ : Span12Mux_h
    port map (
            O => \N__25438\,
            I => \N__25396\
        );

    \I__5174\ : Span4Mux_h
    port map (
            O => \N__25431\,
            I => \N__25391\
        );

    \I__5173\ : Span4Mux_h
    port map (
            O => \N__25428\,
            I => \N__25391\
        );

    \I__5172\ : Span4Mux_h
    port map (
            O => \N__25425\,
            I => \N__25382\
        );

    \I__5171\ : Span4Mux_v
    port map (
            O => \N__25420\,
            I => \N__25382\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__25415\,
            I => \N__25382\
        );

    \I__5169\ : Span4Mux_v
    port map (
            O => \N__25406\,
            I => \N__25382\
        );

    \I__5168\ : CascadeMux
    port map (
            O => \N__25405\,
            I => \N__25379\
        );

    \I__5167\ : CascadeMux
    port map (
            O => \N__25404\,
            I => \N__25375\
        );

    \I__5166\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \N__25371\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__25402\,
            I => \N__25367\
        );

    \I__5164\ : CascadeMux
    port map (
            O => \N__25401\,
            I => \N__25363\
        );

    \I__5163\ : CascadeMux
    port map (
            O => \N__25400\,
            I => \N__25359\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__25399\,
            I => \N__25356\
        );

    \I__5161\ : Span12Mux_v
    port map (
            O => \N__25396\,
            I => \N__25353\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__25391\,
            I => \N__25350\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__25382\,
            I => \N__25347\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25332\
        );

    \I__5157\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25332\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25332\
        );

    \I__5155\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25332\
        );

    \I__5154\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25332\
        );

    \I__5153\ : InMux
    port map (
            O => \N__25370\,
            I => \N__25332\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25332\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25321\
        );

    \I__5150\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25321\
        );

    \I__5149\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25321\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25359\,
            I => \N__25321\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25321\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__25353\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5145\ : Odrv4
    port map (
            O => \N__25350\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5144\ : Odrv4
    port map (
            O => \N__25347\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__25332\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__25321\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25310\,
            I => \M_this_data_count_q_cry_11\
        );

    \I__5140\ : InMux
    port map (
            O => \N__25307\,
            I => \M_this_data_count_q_cry_12\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__5138\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25297\
        );

    \I__5137\ : CascadeMux
    port map (
            O => \N__25300\,
            I => \N__25293\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__25297\,
            I => \N__25288\
        );

    \I__5135\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25285\
        );

    \I__5134\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25278\
        );

    \I__5133\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25278\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25278\
        );

    \I__5131\ : Span4Mux_v
    port map (
            O => \N__25288\,
            I => \N__25275\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__25285\,
            I => \N__25270\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__25278\,
            I => \N__25270\
        );

    \I__5128\ : Span4Mux_v
    port map (
            O => \N__25275\,
            I => \N__25267\
        );

    \I__5127\ : Span4Mux_v
    port map (
            O => \N__25270\,
            I => \N__25264\
        );

    \I__5126\ : Sp12to4
    port map (
            O => \N__25267\,
            I => \N__25259\
        );

    \I__5125\ : Sp12to4
    port map (
            O => \N__25264\,
            I => \N__25259\
        );

    \I__5124\ : Span12Mux_h
    port map (
            O => \N__25259\,
            I => \N__25256\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__25256\,
            I => port_enb_c
        );

    \I__5122\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25250\,
            I => \N__25243\
        );

    \I__5120\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25236\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25248\,
            I => \N__25236\
        );

    \I__5118\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25236\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25233\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__25243\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__25236\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__25233\,
            I => \M_this_delay_clk_out_0\
        );

    \I__5113\ : InMux
    port map (
            O => \N__25226\,
            I => \N__25223\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__5111\ : Odrv4
    port map (
            O => \N__25220\,
            I => \M_this_data_count_q_s_8\
        );

    \I__5110\ : CascadeMux
    port map (
            O => \N__25217\,
            I => \N__25213\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__25216\,
            I => \N__25206\
        );

    \I__5108\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25201\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25201\
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__25211\,
            I => \N__25195\
        );

    \I__5105\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25190\
        );

    \I__5104\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25190\
        );

    \I__5103\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25187\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25184\
        );

    \I__5101\ : InMux
    port map (
            O => \N__25200\,
            I => \N__25179\
        );

    \I__5100\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25179\
        );

    \I__5099\ : CascadeMux
    port map (
            O => \N__25198\,
            I => \N__25176\
        );

    \I__5098\ : InMux
    port map (
            O => \N__25195\,
            I => \N__25173\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__25190\,
            I => \N__25166\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25166\
        );

    \I__5095\ : Span4Mux_h
    port map (
            O => \N__25184\,
            I => \N__25166\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__25179\,
            I => \N__25163\
        );

    \I__5093\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25160\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__25173\,
            I => \N__25157\
        );

    \I__5091\ : Span4Mux_v
    port map (
            O => \N__25166\,
            I => \N__25154\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__25163\,
            I => \N__25149\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__25160\,
            I => \N__25149\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__25157\,
            I => \N_92\
        );

    \I__5087\ : Odrv4
    port map (
            O => \N__25154\,
            I => \N_92\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__25149\,
            I => \N_92\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25142\,
            I => \N__25138\
        );

    \I__5084\ : InMux
    port map (
            O => \N__25141\,
            I => \N__25135\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__25138\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__25135\,
            I => \M_this_data_count_qZ0Z_8\
        );

    \I__5081\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25127\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__25121\,
            I => \M_this_data_count_q_cry_0_THRU_CO\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25118\,
            I => \M_this_data_count_q_cry_0\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25115\,
            I => \N__25112\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__25112\,
            I => \N__25109\
        );

    \I__5074\ : Odrv4
    port map (
            O => \N__25109\,
            I => \M_this_data_count_q_cry_1_THRU_CO\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25106\,
            I => \M_this_data_count_q_cry_1\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25100\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25097\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__25097\,
            I => \M_this_data_count_q_cry_2_THRU_CO\
        );

    \I__5069\ : InMux
    port map (
            O => \N__25094\,
            I => \M_this_data_count_q_cry_2\
        );

    \I__5068\ : InMux
    port map (
            O => \N__25091\,
            I => \M_this_data_count_q_cry_3\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25088\,
            I => \M_this_data_count_q_cry_4\
        );

    \I__5066\ : InMux
    port map (
            O => \N__25085\,
            I => \M_this_data_count_q_cry_5\
        );

    \I__5065\ : CascadeMux
    port map (
            O => \N__25082\,
            I => \N__25079\
        );

    \I__5064\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25076\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5062\ : Odrv4
    port map (
            O => \N__25073\,
            I => \M_this_data_count_q_cry_6_THRU_CO\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25070\,
            I => \M_this_data_count_q_cry_6\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25067\,
            I => \bfn_15_20_0_\
        );

    \I__5059\ : CascadeMux
    port map (
            O => \N__25064\,
            I => \N__25061\
        );

    \I__5058\ : CascadeBuf
    port map (
            O => \N__25061\,
            I => \N__25058\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__25058\,
            I => \N__25055\
        );

    \I__5056\ : InMux
    port map (
            O => \N__25055\,
            I => \N__25052\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__5053\ : Sp12to4
    port map (
            O => \N__25046\,
            I => \N__25041\
        );

    \I__5052\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25038\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25035\
        );

    \I__5050\ : Span12Mux_h
    port map (
            O => \N__25041\,
            I => \N__25032\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25038\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__25035\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5047\ : Odrv12
    port map (
            O => \N__25032\,
            I => \M_this_ppu_map_addr_4\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__5045\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25019\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__5043\ : Odrv4
    port map (
            O => \N__25016\,
            I => \this_ppu.M_oam_cache_read_data_15\
        );

    \I__5042\ : InMux
    port map (
            O => \N__25013\,
            I => \this_ppu.offset_x_cry_6\
        );

    \I__5041\ : InMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__25007\,
            I => \this_ppu.offset_x_7\
        );

    \I__5039\ : CascadeMux
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__5038\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24998\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__24998\,
            I => \M_this_scroll_qZ0Z_0\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24992\
        );

    \I__5035\ : InMux
    port map (
            O => \N__24992\,
            I => \N__24989\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__24989\,
            I => \M_this_scroll_qZ0Z_1\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__24986\,
            I => \N__24983\
        );

    \I__5032\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__24980\,
            I => \M_this_scroll_qZ0Z_2\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__24977\,
            I => \N__24974\
        );

    \I__5029\ : InMux
    port map (
            O => \N__24974\,
            I => \N__24971\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__24971\,
            I => \N__24968\
        );

    \I__5027\ : Odrv12
    port map (
            O => \N__24968\,
            I => \M_this_scroll_qZ0Z_3\
        );

    \I__5026\ : CascadeMux
    port map (
            O => \N__24965\,
            I => \N__24962\
        );

    \I__5025\ : InMux
    port map (
            O => \N__24962\,
            I => \N__24959\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__24959\,
            I => \M_this_scroll_qZ0Z_4\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__24956\,
            I => \N__24953\
        );

    \I__5022\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24950\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__24950\,
            I => \M_this_scroll_qZ0Z_5\
        );

    \I__5020\ : CascadeMux
    port map (
            O => \N__24947\,
            I => \N__24944\
        );

    \I__5019\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__24941\,
            I => \M_this_scroll_qZ0Z_6\
        );

    \I__5017\ : InMux
    port map (
            O => \N__24938\,
            I => \N__24935\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__24935\,
            I => \M_this_scroll_qZ0Z_7\
        );

    \I__5015\ : CascadeMux
    port map (
            O => \N__24932\,
            I => \this_vga_signals.M_vcounter_d7lt8_0_cascade_\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__24929\,
            I => \N__24924\
        );

    \I__5013\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24919\
        );

    \I__5012\ : InMux
    port map (
            O => \N__24927\,
            I => \N__24919\
        );

    \I__5011\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24916\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__24919\,
            I => \N__24909\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__24916\,
            I => \N__24906\
        );

    \I__5008\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24901\
        );

    \I__5007\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24901\
        );

    \I__5006\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24896\
        );

    \I__5005\ : InMux
    port map (
            O => \N__24912\,
            I => \N__24896\
        );

    \I__5004\ : Span4Mux_v
    port map (
            O => \N__24909\,
            I => \N__24891\
        );

    \I__5003\ : Span4Mux_h
    port map (
            O => \N__24906\,
            I => \N__24891\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__24901\,
            I => \this_ppu.offset_x\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__24896\,
            I => \this_ppu.offset_x\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__24891\,
            I => \this_ppu.offset_x\
        );

    \I__4999\ : InMux
    port map (
            O => \N__24884\,
            I => \N__24881\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__24881\,
            I => \this_ppu.M_oam_cache_read_data_i_8\
        );

    \I__4997\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24875\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__24875\,
            I => \N__24872\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__24872\,
            I => \N__24869\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__24869\,
            I => \this_ppu.M_oam_cache_read_data_i_9\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__24866\,
            I => \N__24859\
        );

    \I__4992\ : InMux
    port map (
            O => \N__24865\,
            I => \N__24856\
        );

    \I__4991\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24853\
        );

    \I__4990\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24848\
        );

    \I__4989\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24848\
        );

    \I__4988\ : InMux
    port map (
            O => \N__24859\,
            I => \N__24845\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__24856\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__24853\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__24848\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__24845\,
            I => \this_ppu.M_surface_x_qZ0Z_1\
        );

    \I__4983\ : CascadeMux
    port map (
            O => \N__24836\,
            I => \N__24833\
        );

    \I__4982\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24829\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__24832\,
            I => \N__24826\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24822\
        );

    \I__4979\ : InMux
    port map (
            O => \N__24826\,
            I => \N__24819\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \N__24816\
        );

    \I__4977\ : Span4Mux_h
    port map (
            O => \N__24822\,
            I => \N__24809\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__24819\,
            I => \N__24809\
        );

    \I__4975\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24806\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__24815\,
            I => \N__24803\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__24814\,
            I => \N__24798\
        );

    \I__4972\ : Span4Mux_v
    port map (
            O => \N__24809\,
            I => \N__24791\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__24806\,
            I => \N__24791\
        );

    \I__4970\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24788\
        );

    \I__4969\ : CascadeMux
    port map (
            O => \N__24802\,
            I => \N__24785\
        );

    \I__4968\ : CascadeMux
    port map (
            O => \N__24801\,
            I => \N__24781\
        );

    \I__4967\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24777\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__24797\,
            I => \N__24774\
        );

    \I__4965\ : CascadeMux
    port map (
            O => \N__24796\,
            I => \N__24771\
        );

    \I__4964\ : Span4Mux_v
    port map (
            O => \N__24791\,
            I => \N__24765\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24765\
        );

    \I__4962\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24762\
        );

    \I__4961\ : CascadeMux
    port map (
            O => \N__24784\,
            I => \N__24759\
        );

    \I__4960\ : InMux
    port map (
            O => \N__24781\,
            I => \N__24755\
        );

    \I__4959\ : CascadeMux
    port map (
            O => \N__24780\,
            I => \N__24752\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__24777\,
            I => \N__24749\
        );

    \I__4957\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24746\
        );

    \I__4956\ : InMux
    port map (
            O => \N__24771\,
            I => \N__24743\
        );

    \I__4955\ : CascadeMux
    port map (
            O => \N__24770\,
            I => \N__24740\
        );

    \I__4954\ : Span4Mux_h
    port map (
            O => \N__24765\,
            I => \N__24733\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24733\
        );

    \I__4952\ : InMux
    port map (
            O => \N__24759\,
            I => \N__24730\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__24758\,
            I => \N__24727\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__24755\,
            I => \N__24724\
        );

    \I__4949\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24721\
        );

    \I__4948\ : Span4Mux_h
    port map (
            O => \N__24749\,
            I => \N__24718\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24715\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__24743\,
            I => \N__24712\
        );

    \I__4945\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24709\
        );

    \I__4944\ : CascadeMux
    port map (
            O => \N__24739\,
            I => \N__24706\
        );

    \I__4943\ : CascadeMux
    port map (
            O => \N__24738\,
            I => \N__24703\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__24733\,
            I => \N__24698\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__24730\,
            I => \N__24698\
        );

    \I__4940\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24695\
        );

    \I__4939\ : Span4Mux_h
    port map (
            O => \N__24724\,
            I => \N__24691\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24688\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__24718\,
            I => \N__24683\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__24715\,
            I => \N__24683\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__24712\,
            I => \N__24680\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24677\
        );

    \I__4933\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24674\
        );

    \I__4932\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24671\
        );

    \I__4931\ : Span4Mux_h
    port map (
            O => \N__24698\,
            I => \N__24666\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__24695\,
            I => \N__24666\
        );

    \I__4929\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \N__24663\
        );

    \I__4928\ : Span4Mux_h
    port map (
            O => \N__24691\,
            I => \N__24660\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__24688\,
            I => \N__24657\
        );

    \I__4926\ : Span4Mux_v
    port map (
            O => \N__24683\,
            I => \N__24654\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__24680\,
            I => \N__24649\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__24677\,
            I => \N__24649\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24646\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24643\
        );

    \I__4921\ : Span4Mux_v
    port map (
            O => \N__24666\,
            I => \N__24640\
        );

    \I__4920\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24637\
        );

    \I__4919\ : Sp12to4
    port map (
            O => \N__24660\,
            I => \N__24634\
        );

    \I__4918\ : Span4Mux_h
    port map (
            O => \N__24657\,
            I => \N__24631\
        );

    \I__4917\ : Span4Mux_v
    port map (
            O => \N__24654\,
            I => \N__24628\
        );

    \I__4916\ : Span4Mux_h
    port map (
            O => \N__24649\,
            I => \N__24625\
        );

    \I__4915\ : Span12Mux_s10_h
    port map (
            O => \N__24646\,
            I => \N__24622\
        );

    \I__4914\ : Span12Mux_s9_h
    port map (
            O => \N__24643\,
            I => \N__24619\
        );

    \I__4913\ : Sp12to4
    port map (
            O => \N__24640\,
            I => \N__24614\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24614\
        );

    \I__4911\ : Span12Mux_v
    port map (
            O => \N__24634\,
            I => \N__24609\
        );

    \I__4910\ : Sp12to4
    port map (
            O => \N__24631\,
            I => \N__24609\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__24628\,
            I => \N__24604\
        );

    \I__4908\ : Span4Mux_v
    port map (
            O => \N__24625\,
            I => \N__24604\
        );

    \I__4907\ : Span12Mux_v
    port map (
            O => \N__24622\,
            I => \N__24597\
        );

    \I__4906\ : Span12Mux_v
    port map (
            O => \N__24619\,
            I => \N__24597\
        );

    \I__4905\ : Span12Mux_s10_h
    port map (
            O => \N__24614\,
            I => \N__24597\
        );

    \I__4904\ : Odrv12
    port map (
            O => \N__24609\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__24604\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__4902\ : Odrv12
    port map (
            O => \N__24597\,
            I => \M_this_ppu_spr_addr_1\
        );

    \I__4901\ : InMux
    port map (
            O => \N__24590\,
            I => \this_ppu.offset_x_cry_0\
        );

    \I__4900\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24584\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__24584\,
            I => \N__24581\
        );

    \I__4898\ : Odrv12
    port map (
            O => \N__24581\,
            I => \this_ppu.M_oam_cache_read_data_i_10\
        );

    \I__4897\ : CascadeMux
    port map (
            O => \N__24578\,
            I => \N__24575\
        );

    \I__4896\ : InMux
    port map (
            O => \N__24575\,
            I => \N__24568\
        );

    \I__4895\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24565\
        );

    \I__4894\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24558\
        );

    \I__4893\ : InMux
    port map (
            O => \N__24572\,
            I => \N__24558\
        );

    \I__4892\ : InMux
    port map (
            O => \N__24571\,
            I => \N__24558\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__24568\,
            I => \N__24555\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__24565\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__24558\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__24555\,
            I => \this_ppu.M_surface_x_qZ0Z_2\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__4886\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24541\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__24544\,
            I => \N__24538\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__24541\,
            I => \N__24533\
        );

    \I__4883\ : InMux
    port map (
            O => \N__24538\,
            I => \N__24530\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__24537\,
            I => \N__24527\
        );

    \I__4881\ : CascadeMux
    port map (
            O => \N__24536\,
            I => \N__24522\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__24533\,
            I => \N__24517\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__24530\,
            I => \N__24517\
        );

    \I__4878\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24514\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__24526\,
            I => \N__24511\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__24525\,
            I => \N__24507\
        );

    \I__4875\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24503\
        );

    \I__4874\ : Span4Mux_h
    port map (
            O => \N__24517\,
            I => \N__24496\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__24514\,
            I => \N__24496\
        );

    \I__4872\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24493\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__24510\,
            I => \N__24490\
        );

    \I__4870\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24487\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__24506\,
            I => \N__24484\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__24503\,
            I => \N__24477\
        );

    \I__4867\ : CascadeMux
    port map (
            O => \N__24502\,
            I => \N__24474\
        );

    \I__4866\ : CascadeMux
    port map (
            O => \N__24501\,
            I => \N__24471\
        );

    \I__4865\ : Span4Mux_v
    port map (
            O => \N__24496\,
            I => \N__24466\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24466\
        );

    \I__4863\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24463\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__24487\,
            I => \N__24459\
        );

    \I__4861\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24456\
        );

    \I__4860\ : CascadeMux
    port map (
            O => \N__24483\,
            I => \N__24453\
        );

    \I__4859\ : CascadeMux
    port map (
            O => \N__24482\,
            I => \N__24450\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__24481\,
            I => \N__24447\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__24480\,
            I => \N__24444\
        );

    \I__4856\ : Span4Mux_s2_v
    port map (
            O => \N__24477\,
            I => \N__24440\
        );

    \I__4855\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24437\
        );

    \I__4854\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24434\
        );

    \I__4853\ : Span4Mux_h
    port map (
            O => \N__24466\,
            I => \N__24429\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24429\
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__24462\,
            I => \N__24426\
        );

    \I__4850\ : Span4Mux_s0_v
    port map (
            O => \N__24459\,
            I => \N__24423\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24420\
        );

    \I__4848\ : InMux
    port map (
            O => \N__24453\,
            I => \N__24417\
        );

    \I__4847\ : InMux
    port map (
            O => \N__24450\,
            I => \N__24414\
        );

    \I__4846\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24411\
        );

    \I__4845\ : InMux
    port map (
            O => \N__24444\,
            I => \N__24408\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__24443\,
            I => \N__24405\
        );

    \I__4843\ : Sp12to4
    port map (
            O => \N__24440\,
            I => \N__24400\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24400\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24397\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__24429\,
            I => \N__24394\
        );

    \I__4839\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24391\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__24423\,
            I => \N__24384\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__24420\,
            I => \N__24384\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__24417\,
            I => \N__24384\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24381\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24378\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__24408\,
            I => \N__24375\
        );

    \I__4832\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24372\
        );

    \I__4831\ : Span12Mux_h
    port map (
            O => \N__24400\,
            I => \N__24367\
        );

    \I__4830\ : Span12Mux_h
    port map (
            O => \N__24397\,
            I => \N__24367\
        );

    \I__4829\ : Sp12to4
    port map (
            O => \N__24394\,
            I => \N__24362\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__24391\,
            I => \N__24362\
        );

    \I__4827\ : Sp12to4
    port map (
            O => \N__24384\,
            I => \N__24359\
        );

    \I__4826\ : Sp12to4
    port map (
            O => \N__24381\,
            I => \N__24352\
        );

    \I__4825\ : Sp12to4
    port map (
            O => \N__24378\,
            I => \N__24352\
        );

    \I__4824\ : Sp12to4
    port map (
            O => \N__24375\,
            I => \N__24352\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24372\,
            I => \N__24349\
        );

    \I__4822\ : Span12Mux_v
    port map (
            O => \N__24367\,
            I => \N__24344\
        );

    \I__4821\ : Span12Mux_h
    port map (
            O => \N__24362\,
            I => \N__24344\
        );

    \I__4820\ : Span12Mux_v
    port map (
            O => \N__24359\,
            I => \N__24337\
        );

    \I__4819\ : Span12Mux_v
    port map (
            O => \N__24352\,
            I => \N__24337\
        );

    \I__4818\ : Span12Mux_s11_h
    port map (
            O => \N__24349\,
            I => \N__24337\
        );

    \I__4817\ : Odrv12
    port map (
            O => \N__24344\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__4816\ : Odrv12
    port map (
            O => \N__24337\,
            I => \M_this_ppu_spr_addr_2\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24332\,
            I => \this_ppu.offset_x_cry_1\
        );

    \I__4814\ : CascadeMux
    port map (
            O => \N__24329\,
            I => \N__24325\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__24328\,
            I => \N__24322\
        );

    \I__4812\ : CascadeBuf
    port map (
            O => \N__24325\,
            I => \N__24319\
        );

    \I__4811\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24316\
        );

    \I__4810\ : CascadeMux
    port map (
            O => \N__24319\,
            I => \N__24313\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__24316\,
            I => \N__24310\
        );

    \I__4808\ : InMux
    port map (
            O => \N__24313\,
            I => \N__24307\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__24310\,
            I => \N__24300\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24307\,
            I => \N__24297\
        );

    \I__4805\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24292\
        );

    \I__4804\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24292\
        );

    \I__4803\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24287\
        );

    \I__4802\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24287\
        );

    \I__4801\ : Sp12to4
    port map (
            O => \N__24300\,
            I => \N__24282\
        );

    \I__4800\ : Span12Mux_v
    port map (
            O => \N__24297\,
            I => \N__24282\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__24292\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__24287\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4797\ : Odrv12
    port map (
            O => \N__24282\,
            I => \M_this_ppu_map_addr_0\
        );

    \I__4796\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24272\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__24272\,
            I => \this_ppu.offset_x_3\
        );

    \I__4794\ : InMux
    port map (
            O => \N__24269\,
            I => \this_ppu.offset_x_cry_2\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__24266\,
            I => \N__24263\
        );

    \I__4792\ : CascadeBuf
    port map (
            O => \N__24263\,
            I => \N__24260\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__24260\,
            I => \N__24257\
        );

    \I__4790\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24254\
        );

    \I__4789\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24249\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__24253\,
            I => \N__24246\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__24252\,
            I => \N__24240\
        );

    \I__4786\ : Sp12to4
    port map (
            O => \N__24249\,
            I => \N__24237\
        );

    \I__4785\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24234\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24231\
        );

    \I__4783\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24226\
        );

    \I__4782\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24226\
        );

    \I__4781\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24223\
        );

    \I__4780\ : Span12Mux_v
    port map (
            O => \N__24237\,
            I => \N__24220\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__24234\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__24231\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24226\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__24223\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4775\ : Odrv12
    port map (
            O => \N__24220\,
            I => \M_this_ppu_map_addr_1\
        );

    \I__4774\ : InMux
    port map (
            O => \N__24209\,
            I => \N__24206\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__24206\,
            I => \this_ppu.offset_x_4\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24203\,
            I => \this_ppu.offset_x_cry_3\
        );

    \I__4771\ : InMux
    port map (
            O => \N__24200\,
            I => \N__24197\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__24197\,
            I => \N__24194\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__24191\,
            I => \this_ppu.M_oam_cache_read_data_i_13\
        );

    \I__4767\ : CascadeMux
    port map (
            O => \N__24188\,
            I => \N__24185\
        );

    \I__4766\ : CascadeBuf
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__24182\,
            I => \N__24178\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__24181\,
            I => \N__24175\
        );

    \I__4763\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24172\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24169\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__24172\,
            I => \N__24166\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__24169\,
            I => \N__24160\
        );

    \I__4759\ : Span12Mux_s7_h
    port map (
            O => \N__24166\,
            I => \N__24157\
        );

    \I__4758\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24154\
        );

    \I__4757\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24151\
        );

    \I__4756\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24148\
        );

    \I__4755\ : Span4Mux_h
    port map (
            O => \N__24160\,
            I => \N__24145\
        );

    \I__4754\ : Span12Mux_h
    port map (
            O => \N__24157\,
            I => \N__24142\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__24154\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__24151\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__24148\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4750\ : Odrv4
    port map (
            O => \N__24145\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4749\ : Odrv12
    port map (
            O => \N__24142\,
            I => \M_this_ppu_map_addr_2\
        );

    \I__4748\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24128\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__24128\,
            I => \this_ppu.offset_x_5\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24125\,
            I => \this_ppu.offset_x_cry_4\
        );

    \I__4745\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24119\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__24119\,
            I => \N__24116\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__24116\,
            I => \N__24113\
        );

    \I__4742\ : Odrv4
    port map (
            O => \N__24113\,
            I => \this_ppu.M_oam_cache_read_data_i_14\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__24110\,
            I => \N__24107\
        );

    \I__4740\ : CascadeBuf
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__24104\,
            I => \N__24100\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__24103\,
            I => \N__24097\
        );

    \I__4737\ : InMux
    port map (
            O => \N__24100\,
            I => \N__24094\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24090\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24087\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__24093\,
            I => \N__24083\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__24090\,
            I => \N__24080\
        );

    \I__4732\ : Span12Mux_s7_v
    port map (
            O => \N__24087\,
            I => \N__24077\
        );

    \I__4731\ : InMux
    port map (
            O => \N__24086\,
            I => \N__24072\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24083\,
            I => \N__24072\
        );

    \I__4729\ : Span4Mux_h
    port map (
            O => \N__24080\,
            I => \N__24069\
        );

    \I__4728\ : Span12Mux_h
    port map (
            O => \N__24077\,
            I => \N__24066\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24072\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4726\ : Odrv4
    port map (
            O => \N__24069\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4725\ : Odrv12
    port map (
            O => \N__24066\,
            I => \M_this_ppu_map_addr_3\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24059\,
            I => \N__24056\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__24056\,
            I => \this_ppu.offset_x_6\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24053\,
            I => \this_ppu.offset_x_cry_5\
        );

    \I__4721\ : InMux
    port map (
            O => \N__24050\,
            I => \N__24046\
        );

    \I__4720\ : CascadeMux
    port map (
            O => \N__24049\,
            I => \N__24043\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__24046\,
            I => \N__24040\
        );

    \I__4718\ : InMux
    port map (
            O => \N__24043\,
            I => \N__24037\
        );

    \I__4717\ : Span4Mux_v
    port map (
            O => \N__24040\,
            I => \N__24033\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__24037\,
            I => \N__24030\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24036\,
            I => \N__24027\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__24033\,
            I => \N__24022\
        );

    \I__4713\ : Span4Mux_v
    port map (
            O => \N__24030\,
            I => \N__24022\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__24027\,
            I => \M_this_ctrl_flags_qZ0Z_6\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__24022\,
            I => \M_this_ctrl_flags_qZ0Z_6\
        );

    \I__4710\ : InMux
    port map (
            O => \N__24017\,
            I => \N__24014\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__24014\,
            I => \N__24011\
        );

    \I__4708\ : Span12Mux_v
    port map (
            O => \N__24011\,
            I => \N__24008\
        );

    \I__4707\ : Odrv12
    port map (
            O => \N__24008\,
            I => \M_this_oam_ram_read_data_13\
        );

    \I__4706\ : CEMux
    port map (
            O => \N__24005\,
            I => \N__24002\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23984\
        );

    \I__4704\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23968\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23959\
        );

    \I__4702\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23959\
        );

    \I__4701\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23959\
        );

    \I__4700\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23959\
        );

    \I__4699\ : InMux
    port map (
            O => \N__23996\,
            I => \N__23956\
        );

    \I__4698\ : InMux
    port map (
            O => \N__23995\,
            I => \N__23952\
        );

    \I__4697\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23935\
        );

    \I__4696\ : InMux
    port map (
            O => \N__23993\,
            I => \N__23935\
        );

    \I__4695\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23935\
        );

    \I__4694\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23935\
        );

    \I__4693\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23935\
        );

    \I__4692\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23935\
        );

    \I__4691\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23935\
        );

    \I__4690\ : InMux
    port map (
            O => \N__23987\,
            I => \N__23932\
        );

    \I__4689\ : Span4Mux_v
    port map (
            O => \N__23984\,
            I => \N__23929\
        );

    \I__4688\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23924\
        );

    \I__4687\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23924\
        );

    \I__4686\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23913\
        );

    \I__4685\ : InMux
    port map (
            O => \N__23980\,
            I => \N__23913\
        );

    \I__4684\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23913\
        );

    \I__4683\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23913\
        );

    \I__4682\ : InMux
    port map (
            O => \N__23977\,
            I => \N__23913\
        );

    \I__4681\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23904\
        );

    \I__4680\ : InMux
    port map (
            O => \N__23975\,
            I => \N__23904\
        );

    \I__4679\ : InMux
    port map (
            O => \N__23974\,
            I => \N__23904\
        );

    \I__4678\ : InMux
    port map (
            O => \N__23973\,
            I => \N__23904\
        );

    \I__4677\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23899\
        );

    \I__4676\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23899\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__23968\,
            I => \N__23894\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23894\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__23956\,
            I => \N__23891\
        );

    \I__4672\ : InMux
    port map (
            O => \N__23955\,
            I => \N__23888\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23879\
        );

    \I__4670\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23876\
        );

    \I__4669\ : CEMux
    port map (
            O => \N__23950\,
            I => \N__23873\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23870\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__23932\,
            I => \N__23867\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__23929\,
            I => \N__23860\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__23924\,
            I => \N__23860\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__23913\,
            I => \N__23860\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__23904\,
            I => \N__23855\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__23899\,
            I => \N__23855\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__23894\,
            I => \N__23850\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__23891\,
            I => \N__23850\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__23888\,
            I => \N__23846\
        );

    \I__4658\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23839\
        );

    \I__4657\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23839\
        );

    \I__4656\ : InMux
    port map (
            O => \N__23885\,
            I => \N__23839\
        );

    \I__4655\ : InMux
    port map (
            O => \N__23884\,
            I => \N__23832\
        );

    \I__4654\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23832\
        );

    \I__4653\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23832\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__23879\,
            I => \N__23827\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23827\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__23873\,
            I => \N__23824\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__23870\,
            I => \N__23817\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__23867\,
            I => \N__23817\
        );

    \I__4647\ : Span4Mux_v
    port map (
            O => \N__23860\,
            I => \N__23817\
        );

    \I__4646\ : Span12Mux_s6_v
    port map (
            O => \N__23855\,
            I => \N__23814\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__23850\,
            I => \N__23811\
        );

    \I__4644\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23808\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__23846\,
            I => \N__23805\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23798\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__23832\,
            I => \N__23798\
        );

    \I__4640\ : Span4Mux_h
    port map (
            O => \N__23827\,
            I => \N__23798\
        );

    \I__4639\ : Odrv12
    port map (
            O => \N__23824\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__23817\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__23814\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4636\ : Odrv4
    port map (
            O => \N__23811\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__23808\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__23805\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__23798\,
            I => \this_ppu.M_state_qZ0Z_3\
        );

    \I__4632\ : InMux
    port map (
            O => \N__23783\,
            I => \N__23780\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23777\
        );

    \I__4630\ : Span4Mux_v
    port map (
            O => \N__23777\,
            I => \N__23774\
        );

    \I__4629\ : Span4Mux_v
    port map (
            O => \N__23774\,
            I => \N__23771\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__23771\,
            I => \N__23768\
        );

    \I__4627\ : Odrv4
    port map (
            O => \N__23768\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_13\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__23765\,
            I => \N__23760\
        );

    \I__4625\ : InMux
    port map (
            O => \N__23764\,
            I => \N__23752\
        );

    \I__4624\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23752\
        );

    \I__4623\ : InMux
    port map (
            O => \N__23760\,
            I => \N__23749\
        );

    \I__4622\ : InMux
    port map (
            O => \N__23759\,
            I => \N__23746\
        );

    \I__4621\ : InMux
    port map (
            O => \N__23758\,
            I => \N__23743\
        );

    \I__4620\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23740\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__23752\,
            I => \N__23737\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__23749\,
            I => \N__23734\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__23746\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__23743\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__23740\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4614\ : Odrv4
    port map (
            O => \N__23737\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4613\ : Odrv4
    port map (
            O => \N__23734\,
            I => \M_this_oam_address_qZ0Z_1\
        );

    \I__4612\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23716\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23713\
        );

    \I__4610\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23710\
        );

    \I__4609\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23705\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23719\,
            I => \N__23705\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23699\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__23713\,
            I => \N__23699\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__23710\,
            I => \N__23694\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23694\
        );

    \I__4603\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23690\
        );

    \I__4602\ : Span4Mux_h
    port map (
            O => \N__23699\,
            I => \N__23687\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__23694\,
            I => \N__23684\
        );

    \I__4600\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23681\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__23690\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__23687\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__23684\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__23681\,
            I => \M_this_oam_address_qZ0Z_0\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__23672\,
            I => \N__23668\
        );

    \I__4594\ : CascadeMux
    port map (
            O => \N__23671\,
            I => \N__23664\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23659\
        );

    \I__4592\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23655\
        );

    \I__4591\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23652\
        );

    \I__4590\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23647\
        );

    \I__4589\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23647\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__23659\,
            I => \N__23644\
        );

    \I__4587\ : InMux
    port map (
            O => \N__23658\,
            I => \N__23641\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__23655\,
            I => \N__23634\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__23652\,
            I => \N__23634\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23634\
        );

    \I__4583\ : Span4Mux_v
    port map (
            O => \N__23644\,
            I => \N__23631\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__23641\,
            I => \N__23626\
        );

    \I__4581\ : Span4Mux_v
    port map (
            O => \N__23634\,
            I => \N__23626\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__23631\,
            I => \N_222_0\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__23626\,
            I => \N_222_0\
        );

    \I__4578\ : CEMux
    port map (
            O => \N__23621\,
            I => \N__23616\
        );

    \I__4577\ : CEMux
    port map (
            O => \N__23620\,
            I => \N__23613\
        );

    \I__4576\ : CEMux
    port map (
            O => \N__23619\,
            I => \N__23610\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__23616\,
            I => \N__23607\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23603\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__23610\,
            I => \N__23600\
        );

    \I__4572\ : Span4Mux_v
    port map (
            O => \N__23607\,
            I => \N__23597\
        );

    \I__4571\ : CEMux
    port map (
            O => \N__23606\,
            I => \N__23594\
        );

    \I__4570\ : Span4Mux_v
    port map (
            O => \N__23603\,
            I => \N__23589\
        );

    \I__4569\ : Span4Mux_v
    port map (
            O => \N__23600\,
            I => \N__23589\
        );

    \I__4568\ : Span4Mux_h
    port map (
            O => \N__23597\,
            I => \N__23584\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__23594\,
            I => \N__23584\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__23589\,
            I => \N__23581\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__23584\,
            I => \N__23578\
        );

    \I__4564\ : Odrv4
    port map (
            O => \N__23581\,
            I => \N_1248_0\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__23578\,
            I => \N_1248_0\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23570\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__23570\,
            I => \this_reset_cond.M_stage_qZ0Z_2\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__23567\,
            I => \M_this_spr_ram_write_en_0_i_1_0_cascade_\
        );

    \I__4559\ : CEMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23558\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__23558\,
            I => \N__23554\
        );

    \I__4556\ : CEMux
    port map (
            O => \N__23557\,
            I => \N__23551\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__23551\,
            I => \N__23545\
        );

    \I__4553\ : Sp12to4
    port map (
            O => \N__23548\,
            I => \N__23542\
        );

    \I__4552\ : Sp12to4
    port map (
            O => \N__23545\,
            I => \N__23539\
        );

    \I__4551\ : Span12Mux_v
    port map (
            O => \N__23542\,
            I => \N__23534\
        );

    \I__4550\ : Span12Mux_v
    port map (
            O => \N__23539\,
            I => \N__23534\
        );

    \I__4549\ : Odrv12
    port map (
            O => \N__23534\,
            I => \this_spr_ram.mem_WE_2\
        );

    \I__4548\ : InMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23525\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__23525\,
            I => \N__23522\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__23522\,
            I => \this_vga_signals.M_vcounter_d7lt8_0\
        );

    \I__4544\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23516\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__23516\,
            I => \N__23513\
        );

    \I__4542\ : Span4Mux_h
    port map (
            O => \N__23513\,
            I => \N__23510\
        );

    \I__4541\ : Span4Mux_h
    port map (
            O => \N__23510\,
            I => \N__23507\
        );

    \I__4540\ : Span4Mux_h
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__4539\ : Odrv4
    port map (
            O => \N__23504\,
            I => \this_delay_clk.M_pipe_qZ0Z_3\
        );

    \I__4538\ : CEMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23495\
        );

    \I__4536\ : Span4Mux_h
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__23492\,
            I => \N_1256_0\
        );

    \I__4534\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23486\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__4532\ : Span4Mux_h
    port map (
            O => \N__23483\,
            I => \N__23479\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23476\
        );

    \I__4530\ : Sp12to4
    port map (
            O => \N__23479\,
            I => \N__23473\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__23476\,
            I => \N__23470\
        );

    \I__4528\ : Span12Mux_v
    port map (
            O => \N__23473\,
            I => \N__23467\
        );

    \I__4527\ : Span12Mux_v
    port map (
            O => \N__23470\,
            I => \N__23464\
        );

    \I__4526\ : Odrv12
    port map (
            O => \N__23467\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__4525\ : Odrv12
    port map (
            O => \N__23464\,
            I => \M_this_oam_ram_read_data_16\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23456\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__23456\,
            I => \N__23453\
        );

    \I__4522\ : Span4Mux_v
    port map (
            O => \N__23453\,
            I => \N__23450\
        );

    \I__4521\ : Span4Mux_h
    port map (
            O => \N__23450\,
            I => \N__23447\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__23447\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_16\
        );

    \I__4519\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23441\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23438\
        );

    \I__4517\ : Span4Mux_v
    port map (
            O => \N__23438\,
            I => \N__23434\
        );

    \I__4516\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23431\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__23434\,
            I => \N__23426\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23426\
        );

    \I__4513\ : Sp12to4
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__4512\ : Span12Mux_v
    port map (
            O => \N__23423\,
            I => \N__23420\
        );

    \I__4511\ : Odrv12
    port map (
            O => \N__23420\,
            I => \M_this_oam_ram_read_data_17\
        );

    \I__4510\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23414\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23411\
        );

    \I__4508\ : Span4Mux_v
    port map (
            O => \N__23411\,
            I => \N__23408\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__23408\,
            I => \N__23405\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__23405\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_17\
        );

    \I__4505\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23399\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__23399\,
            I => \N__23395\
        );

    \I__4503\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23392\
        );

    \I__4502\ : Span4Mux_h
    port map (
            O => \N__23395\,
            I => \N__23389\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__23392\,
            I => \N__23386\
        );

    \I__4500\ : Sp12to4
    port map (
            O => \N__23389\,
            I => \N__23383\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__23386\,
            I => \N__23380\
        );

    \I__4498\ : Span12Mux_v
    port map (
            O => \N__23383\,
            I => \N__23377\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__23380\,
            I => \N__23374\
        );

    \I__4496\ : Odrv12
    port map (
            O => \N__23377\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__23374\,
            I => \M_this_oam_ram_read_data_18\
        );

    \I__4494\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23366\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N__23363\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__23363\,
            I => \N__23360\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__23360\,
            I => \N__23357\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__23357\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_18\
        );

    \I__4489\ : InMux
    port map (
            O => \N__23354\,
            I => \N__23351\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__23351\,
            I => \N__23348\
        );

    \I__4487\ : Span4Mux_h
    port map (
            O => \N__23348\,
            I => \N__23345\
        );

    \I__4486\ : Sp12to4
    port map (
            O => \N__23345\,
            I => \N__23342\
        );

    \I__4485\ : Span12Mux_v
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__4484\ : Odrv12
    port map (
            O => \N__23339\,
            I => \M_this_oam_ram_read_data_27\
        );

    \I__4483\ : InMux
    port map (
            O => \N__23336\,
            I => \N__23333\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23333\,
            I => \N__23330\
        );

    \I__4481\ : Odrv12
    port map (
            O => \N__23330\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_27\
        );

    \I__4480\ : InMux
    port map (
            O => \N__23327\,
            I => \this_ppu.un1_M_surface_y_d_cry_5\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__23324\,
            I => \N__23321\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23321\,
            I => \N__23317\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__23320\,
            I => \N__23314\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__23317\,
            I => \N__23311\
        );

    \I__4475\ : InMux
    port map (
            O => \N__23314\,
            I => \N__23308\
        );

    \I__4474\ : Odrv12
    port map (
            O => \N__23311\,
            I => \this_ppu.M_screen_y_qZ0Z_7\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__23308\,
            I => \this_ppu.M_screen_y_qZ0Z_7\
        );

    \I__4472\ : InMux
    port map (
            O => \N__23303\,
            I => \bfn_14_19_0_\
        );

    \I__4471\ : CascadeMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__4470\ : CascadeBuf
    port map (
            O => \N__23297\,
            I => \N__23293\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23296\,
            I => \N__23290\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__23293\,
            I => \N__23287\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__23290\,
            I => \N__23284\
        );

    \I__4466\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__23284\,
            I => \N__23278\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23275\
        );

    \I__4463\ : Span4Mux_h
    port map (
            O => \N__23278\,
            I => \N__23272\
        );

    \I__4462\ : Span12Mux_h
    port map (
            O => \N__23275\,
            I => \N__23269\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__23272\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4460\ : Odrv12
    port map (
            O => \N__23269\,
            I => \M_this_ppu_map_addr_9\
        );

    \I__4459\ : CascadeMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__4458\ : InMux
    port map (
            O => \N__23261\,
            I => \N__23258\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23250\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__23257\,
            I => \N__23247\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23242\
        );

    \I__4454\ : InMux
    port map (
            O => \N__23255\,
            I => \N__23242\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23254\,
            I => \N__23236\
        );

    \I__4452\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23236\
        );

    \I__4451\ : Span12Mux_v
    port map (
            O => \N__23250\,
            I => \N__23233\
        );

    \I__4450\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23230\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23227\
        );

    \I__4448\ : InMux
    port map (
            O => \N__23241\,
            I => \N__23224\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23221\
        );

    \I__4446\ : Odrv12
    port map (
            O => \N__23233\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__23230\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__23227\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__23224\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__23221\,
            I => \M_this_ppu_vram_addr_7\
        );

    \I__4441\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23204\
        );

    \I__4440\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23201\
        );

    \I__4439\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23196\
        );

    \I__4438\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23196\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__23204\,
            I => \N__23193\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__23201\,
            I => \N__23190\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__23196\,
            I => \this_ppu.M_screen_y_qZ0Z_1\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__23193\,
            I => \this_ppu.M_screen_y_qZ0Z_1\
        );

    \I__4433\ : Odrv12
    port map (
            O => \N__23190\,
            I => \this_ppu.M_screen_y_qZ0Z_1\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__23183\,
            I => \N__23172\
        );

    \I__4431\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23168\
        );

    \I__4430\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23159\
        );

    \I__4429\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23159\
        );

    \I__4428\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23159\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23159\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23177\,
            I => \N__23151\
        );

    \I__4425\ : InMux
    port map (
            O => \N__23176\,
            I => \N__23151\
        );

    \I__4424\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23151\
        );

    \I__4423\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23148\
        );

    \I__4422\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23145\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23133\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__23159\,
            I => \N__23133\
        );

    \I__4419\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23130\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__23151\,
            I => \N__23123\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__23148\,
            I => \N__23123\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23123\
        );

    \I__4415\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23114\
        );

    \I__4414\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23114\
        );

    \I__4413\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23114\
        );

    \I__4412\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23114\
        );

    \I__4411\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23107\
        );

    \I__4410\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23107\
        );

    \I__4409\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23107\
        );

    \I__4408\ : Odrv4
    port map (
            O => \N__23133\,
            I => \M_this_ppu_vga_is_drawing\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__23130\,
            I => \M_this_ppu_vga_is_drawing\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__23123\,
            I => \M_this_ppu_vga_is_drawing\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__23114\,
            I => \M_this_ppu_vga_is_drawing\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__23107\,
            I => \M_this_ppu_vga_is_drawing\
        );

    \I__4403\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23091\
        );

    \I__4402\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23087\
        );

    \I__4401\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23084\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__23091\,
            I => \N__23081\
        );

    \I__4399\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23078\
        );

    \I__4398\ : InMux
    port map (
            O => \N__23087\,
            I => \N__23075\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23072\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__23081\,
            I => \N__23067\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__23078\,
            I => \N__23067\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__23075\,
            I => \this_ppu.M_screen_y_qZ0Z_2\
        );

    \I__4393\ : Odrv12
    port map (
            O => \N__23072\,
            I => \this_ppu.M_screen_y_qZ0Z_2\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__23067\,
            I => \this_ppu.M_screen_y_qZ0Z_2\
        );

    \I__4391\ : CEMux
    port map (
            O => \N__23060\,
            I => \N__23055\
        );

    \I__4390\ : CEMux
    port map (
            O => \N__23059\,
            I => \N__23052\
        );

    \I__4389\ : CEMux
    port map (
            O => \N__23058\,
            I => \N__23048\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__23055\,
            I => \N__23045\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23042\
        );

    \I__4386\ : CEMux
    port map (
            O => \N__23051\,
            I => \N__23039\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__23036\
        );

    \I__4384\ : Span4Mux_v
    port map (
            O => \N__23045\,
            I => \N__23029\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__23042\,
            I => \N__23029\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__23039\,
            I => \N__23029\
        );

    \I__4381\ : Span4Mux_h
    port map (
            O => \N__23036\,
            I => \N__23026\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__23029\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__23026\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0\
        );

    \I__4378\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23018\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__23018\,
            I => \N__23015\
        );

    \I__4376\ : Span12Mux_h
    port map (
            O => \N__23015\,
            I => \N__23012\
        );

    \I__4375\ : Odrv12
    port map (
            O => \N__23012\,
            I => \M_this_oam_ram_read_data_12\
        );

    \I__4374\ : InMux
    port map (
            O => \N__23009\,
            I => \N__23006\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__23006\,
            I => \N__23003\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__23003\,
            I => \N__23000\
        );

    \I__4371\ : Span4Mux_h
    port map (
            O => \N__23000\,
            I => \N__22997\
        );

    \I__4370\ : Odrv4
    port map (
            O => \N__22997\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_12\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22990\
        );

    \I__4368\ : CascadeMux
    port map (
            O => \N__22993\,
            I => \N__22984\
        );

    \I__4367\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22979\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__22989\,
            I => \N__22976\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__22988\,
            I => \N__22973\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__22987\,
            I => \N__22968\
        );

    \I__4363\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22964\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__22983\,
            I => \N__22961\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__22982\,
            I => \N__22958\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22954\
        );

    \I__4359\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22951\
        );

    \I__4358\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22948\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__22972\,
            I => \N__22945\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__22971\,
            I => \N__22942\
        );

    \I__4355\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22937\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__22967\,
            I => \N__22934\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__22964\,
            I => \N__22931\
        );

    \I__4352\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22928\
        );

    \I__4351\ : InMux
    port map (
            O => \N__22958\,
            I => \N__22925\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__22957\,
            I => \N__22922\
        );

    \I__4349\ : Span4Mux_s0_v
    port map (
            O => \N__22954\,
            I => \N__22916\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__22951\,
            I => \N__22916\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22913\
        );

    \I__4346\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22910\
        );

    \I__4345\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22907\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__22941\,
            I => \N__22904\
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__22940\,
            I => \N__22901\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__22937\,
            I => \N__22897\
        );

    \I__4341\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22894\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__22931\,
            I => \N__22891\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__22928\,
            I => \N__22888\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22885\
        );

    \I__4337\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22882\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__22921\,
            I => \N__22879\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__22916\,
            I => \N__22872\
        );

    \I__4334\ : Span4Mux_h
    port map (
            O => \N__22913\,
            I => \N__22872\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__22910\,
            I => \N__22872\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__22907\,
            I => \N__22869\
        );

    \I__4331\ : InMux
    port map (
            O => \N__22904\,
            I => \N__22866\
        );

    \I__4330\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22863\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \N__22860\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__22897\,
            I => \N__22856\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__22894\,
            I => \N__22853\
        );

    \I__4326\ : Span4Mux_v
    port map (
            O => \N__22891\,
            I => \N__22848\
        );

    \I__4325\ : Span4Mux_h
    port map (
            O => \N__22888\,
            I => \N__22848\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__22885\,
            I => \N__22845\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__22882\,
            I => \N__22842\
        );

    \I__4322\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22839\
        );

    \I__4321\ : Span4Mux_v
    port map (
            O => \N__22872\,
            I => \N__22832\
        );

    \I__4320\ : Span4Mux_h
    port map (
            O => \N__22869\,
            I => \N__22832\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22832\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22829\
        );

    \I__4317\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22826\
        );

    \I__4316\ : CascadeMux
    port map (
            O => \N__22859\,
            I => \N__22823\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__22856\,
            I => \N__22820\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__22853\,
            I => \N__22817\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__22848\,
            I => \N__22814\
        );

    \I__4312\ : Span4Mux_v
    port map (
            O => \N__22845\,
            I => \N__22809\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__22842\,
            I => \N__22809\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__22839\,
            I => \N__22806\
        );

    \I__4309\ : Span4Mux_v
    port map (
            O => \N__22832\,
            I => \N__22799\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__22829\,
            I => \N__22799\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22799\
        );

    \I__4306\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22796\
        );

    \I__4305\ : Sp12to4
    port map (
            O => \N__22820\,
            I => \N__22793\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__22817\,
            I => \N__22790\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__22814\,
            I => \N__22787\
        );

    \I__4302\ : Span4Mux_h
    port map (
            O => \N__22809\,
            I => \N__22784\
        );

    \I__4301\ : Span12Mux_s10_h
    port map (
            O => \N__22806\,
            I => \N__22781\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__22799\,
            I => \N__22778\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__22796\,
            I => \N__22775\
        );

    \I__4298\ : Span12Mux_s11_v
    port map (
            O => \N__22793\,
            I => \N__22770\
        );

    \I__4297\ : Sp12to4
    port map (
            O => \N__22790\,
            I => \N__22770\
        );

    \I__4296\ : Span4Mux_h
    port map (
            O => \N__22787\,
            I => \N__22765\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__22784\,
            I => \N__22765\
        );

    \I__4294\ : Span12Mux_v
    port map (
            O => \N__22781\,
            I => \N__22758\
        );

    \I__4293\ : Sp12to4
    port map (
            O => \N__22778\,
            I => \N__22758\
        );

    \I__4292\ : Span12Mux_s9_h
    port map (
            O => \N__22775\,
            I => \N__22758\
        );

    \I__4291\ : Odrv12
    port map (
            O => \N__22770\,
            I => \M_this_ppu_spr_addr_8\
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__22765\,
            I => \M_this_ppu_spr_addr_8\
        );

    \I__4289\ : Odrv12
    port map (
            O => \N__22758\,
            I => \M_this_ppu_spr_addr_8\
        );

    \I__4288\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__22748\,
            I => \N__22745\
        );

    \I__4286\ : Odrv4
    port map (
            O => \N__22745\,
            I => \this_ppu.M_screen_y_q_RNICCMV8Z0Z_0\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__22742\,
            I => \N__22738\
        );

    \I__4284\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22734\
        );

    \I__4283\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22731\
        );

    \I__4282\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22728\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22723\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22723\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22720\
        );

    \I__4278\ : Span4Mux_v
    port map (
            O => \N__22723\,
            I => \N__22717\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__22720\,
            I => \N__22714\
        );

    \I__4276\ : Span4Mux_h
    port map (
            O => \N__22717\,
            I => \N__22711\
        );

    \I__4275\ : Odrv4
    port map (
            O => \N__22714\,
            I => \this_ppu.offset_y\
        );

    \I__4274\ : Odrv4
    port map (
            O => \N__22711\,
            I => \this_ppu.offset_y\
        );

    \I__4273\ : InMux
    port map (
            O => \N__22706\,
            I => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\
        );

    \I__4272\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22700\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__22697\,
            I => \this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__22694\,
            I => \N__22690\
        );

    \I__4268\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22687\
        );

    \I__4267\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22684\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__22687\,
            I => \N__22681\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22678\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__22681\,
            I => \N__22673\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__22678\,
            I => \N__22673\
        );

    \I__4262\ : Span4Mux_h
    port map (
            O => \N__22673\,
            I => \N__22670\
        );

    \I__4261\ : Odrv4
    port map (
            O => \N__22670\,
            I => \this_ppu.M_surface_y_qZ0Z_1\
        );

    \I__4260\ : InMux
    port map (
            O => \N__22667\,
            I => \this_ppu.un1_M_surface_y_d_cry_0\
        );

    \I__4259\ : InMux
    port map (
            O => \N__22664\,
            I => \N__22661\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__22661\,
            I => \N__22658\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__22658\,
            I => \N__22655\
        );

    \I__4256\ : Odrv4
    port map (
            O => \N__22655\,
            I => \this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__22652\,
            I => \N__22648\
        );

    \I__4254\ : InMux
    port map (
            O => \N__22651\,
            I => \N__22645\
        );

    \I__4253\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22642\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__22645\,
            I => \N__22639\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__22642\,
            I => \N__22636\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__22639\,
            I => \N__22633\
        );

    \I__4249\ : Span12Mux_h
    port map (
            O => \N__22636\,
            I => \N__22630\
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__22633\,
            I => \this_ppu.M_surface_y_qZ0Z_2\
        );

    \I__4247\ : Odrv12
    port map (
            O => \N__22630\,
            I => \this_ppu.M_surface_y_qZ0Z_2\
        );

    \I__4246\ : InMux
    port map (
            O => \N__22625\,
            I => \this_ppu.un1_M_surface_y_d_cry_1\
        );

    \I__4245\ : InMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__22616\,
            I => \this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__4241\ : CascadeBuf
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__4240\ : CascadeMux
    port map (
            O => \N__22607\,
            I => \N__22603\
        );

    \I__4239\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \N__22600\
        );

    \I__4238\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22597\
        );

    \I__4237\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22594\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__22597\,
            I => \N__22591\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__22594\,
            I => \N__22588\
        );

    \I__4234\ : Span4Mux_v
    port map (
            O => \N__22591\,
            I => \N__22585\
        );

    \I__4233\ : Span4Mux_h
    port map (
            O => \N__22588\,
            I => \N__22582\
        );

    \I__4232\ : Sp12to4
    port map (
            O => \N__22585\,
            I => \N__22579\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__22582\,
            I => \N__22576\
        );

    \I__4230\ : Span12Mux_v
    port map (
            O => \N__22579\,
            I => \N__22573\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__22576\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4228\ : Odrv12
    port map (
            O => \N__22573\,
            I => \M_this_ppu_map_addr_5\
        );

    \I__4227\ : InMux
    port map (
            O => \N__22568\,
            I => \this_ppu.un1_M_surface_y_d_cry_2\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__4224\ : Odrv4
    port map (
            O => \N__22559\,
            I => \this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__22556\,
            I => \N__22552\
        );

    \I__4222\ : CascadeMux
    port map (
            O => \N__22555\,
            I => \N__22549\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__22552\,
            I => \N__22546\
        );

    \I__4220\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22543\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__22546\,
            I => \N__22540\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22537\
        );

    \I__4217\ : InMux
    port map (
            O => \N__22540\,
            I => \N__22534\
        );

    \I__4216\ : Span4Mux_h
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22528\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__22531\,
            I => \N__22525\
        );

    \I__4213\ : Span12Mux_v
    port map (
            O => \N__22528\,
            I => \N__22522\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__22525\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4211\ : Odrv12
    port map (
            O => \N__22522\,
            I => \M_this_ppu_map_addr_6\
        );

    \I__4210\ : InMux
    port map (
            O => \N__22517\,
            I => \this_ppu.un1_M_surface_y_d_cry_3\
        );

    \I__4209\ : InMux
    port map (
            O => \N__22514\,
            I => \N__22511\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__22511\,
            I => \N__22508\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__22508\,
            I => \this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__22505\,
            I => \N__22502\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__22502\,
            I => \N__22499\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__22499\,
            I => \N__22496\
        );

    \I__4203\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22492\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__22495\,
            I => \N__22489\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__22492\,
            I => \N__22486\
        );

    \I__4200\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22483\
        );

    \I__4199\ : Span4Mux_v
    port map (
            O => \N__22486\,
            I => \N__22480\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22477\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__22480\,
            I => \N__22474\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__22477\,
            I => \N__22471\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__22474\,
            I => \N__22468\
        );

    \I__4194\ : Span4Mux_h
    port map (
            O => \N__22471\,
            I => \N__22465\
        );

    \I__4193\ : Sp12to4
    port map (
            O => \N__22468\,
            I => \N__22462\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__22465\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4191\ : Odrv12
    port map (
            O => \N__22462\,
            I => \M_this_ppu_map_addr_7\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22457\,
            I => \this_ppu.un1_M_surface_y_d_cry_4\
        );

    \I__4189\ : InMux
    port map (
            O => \N__22454\,
            I => \N__22451\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__22448\,
            I => \this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6\
        );

    \I__4186\ : CascadeMux
    port map (
            O => \N__22445\,
            I => \N__22442\
        );

    \I__4185\ : CascadeBuf
    port map (
            O => \N__22442\,
            I => \N__22439\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__22439\,
            I => \N__22435\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__22438\,
            I => \N__22432\
        );

    \I__4182\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22429\
        );

    \I__4181\ : InMux
    port map (
            O => \N__22432\,
            I => \N__22426\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22429\,
            I => \N__22423\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22420\
        );

    \I__4178\ : Sp12to4
    port map (
            O => \N__22423\,
            I => \N__22417\
        );

    \I__4177\ : Span4Mux_h
    port map (
            O => \N__22420\,
            I => \N__22414\
        );

    \I__4176\ : Span12Mux_s7_v
    port map (
            O => \N__22417\,
            I => \N__22411\
        );

    \I__4175\ : Span4Mux_h
    port map (
            O => \N__22414\,
            I => \N__22408\
        );

    \I__4174\ : Span12Mux_h
    port map (
            O => \N__22411\,
            I => \N__22405\
        );

    \I__4173\ : Odrv4
    port map (
            O => \N__22408\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__4172\ : Odrv12
    port map (
            O => \N__22405\,
            I => \M_this_ppu_map_addr_8\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__22400\,
            I => \M_this_ppu_vga_is_drawing_cascade_\
        );

    \I__4170\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22393\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__22396\,
            I => \N__22389\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22386\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22382\
        );

    \I__4166\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22379\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__22386\,
            I => \N__22376\
        );

    \I__4164\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22373\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__22382\,
            I => \N__22370\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__22379\,
            I => \this_ppu_M_screen_y_q_5\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__22376\,
            I => \this_ppu_M_screen_y_q_5\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__22373\,
            I => \this_ppu_M_screen_y_q_5\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__22370\,
            I => \this_ppu_M_screen_y_q_5\
        );

    \I__4158\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22358\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__22358\,
            I => \N__22352\
        );

    \I__4156\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22349\
        );

    \I__4155\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22344\
        );

    \I__4154\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22344\
        );

    \I__4153\ : Span4Mux_h
    port map (
            O => \N__22352\,
            I => \N__22339\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22339\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__22344\,
            I => \this_ppu_M_screen_y_q_6\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__22339\,
            I => \this_ppu_M_screen_y_q_6\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22331\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__22331\,
            I => \this_ppu.un1_M_surface_x_q_c1\
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__4146\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__4144\ : Span4Mux_v
    port map (
            O => \N__22319\,
            I => \N__22316\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__22316\,
            I => \M_this_scroll_qZ0Z_9\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22307\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__22307\,
            I => \M_this_scroll_qZ0Z_15\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22301\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__22301\,
            I => \N__22298\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__22298\,
            I => \this_ppu.un1_M_surface_x_q_ac0_11\
        );

    \I__4136\ : InMux
    port map (
            O => \N__22295\,
            I => \N__22292\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__22292\,
            I => \N__22289\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__22289\,
            I => \M_this_scroll_qZ0Z_12\
        );

    \I__4133\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22282\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22285\,
            I => \N__22279\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__22282\,
            I => \this_ppu.un1_M_surface_x_q_c4\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__22279\,
            I => \this_ppu.un1_M_surface_x_q_c4\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__22274\,
            I => \N__22271\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22271\,
            I => \N__22263\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22270\,
            I => \N__22258\
        );

    \I__4126\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22258\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22244\
        );

    \I__4124\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22244\
        );

    \I__4123\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22241\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22263\,
            I => \N__22236\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__22258\,
            I => \N__22236\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22225\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22225\
        );

    \I__4118\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22225\
        );

    \I__4117\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22225\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22225\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22220\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22220\
        );

    \I__4113\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22215\
        );

    \I__4112\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22215\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22210\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__22241\,
            I => \N__22210\
        );

    \I__4109\ : Span4Mux_v
    port map (
            O => \N__22236\,
            I => \N__22207\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__22225\,
            I => \N__22204\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__22220\,
            I => \N__22199\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__22215\,
            I => \N__22199\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__22210\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__22207\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\
        );

    \I__4103\ : Odrv4
    port map (
            O => \N__22204\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__22199\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\
        );

    \I__4101\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__4098\ : Odrv4
    port map (
            O => \N__22181\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_2\
        );

    \I__4097\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22175\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__4095\ : Sp12to4
    port map (
            O => \N__22172\,
            I => \N__22169\
        );

    \I__4094\ : Span12Mux_v
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__4093\ : Odrv12
    port map (
            O => \N__22166\,
            I => \M_this_map_ram_read_data_2\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22163\,
            I => \N__22159\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22156\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22159\,
            I => \this_ppu.un3_M_screen_y_d_0_c6\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__22156\,
            I => \this_ppu.un3_M_screen_y_d_0_c6\
        );

    \I__4088\ : InMux
    port map (
            O => \N__22151\,
            I => \N__22147\
        );

    \I__4087\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22144\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__22147\,
            I => \N__22141\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__22144\,
            I => \this_ppu.un3_M_screen_y_d_0_c4\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__22141\,
            I => \this_ppu.un3_M_screen_y_d_0_c4\
        );

    \I__4083\ : InMux
    port map (
            O => \N__22136\,
            I => \N__22131\
        );

    \I__4082\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22128\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__22134\,
            I => \N__22125\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__22131\,
            I => \N__22120\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__22128\,
            I => \N__22120\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22115\
        );

    \I__4077\ : Span4Mux_v
    port map (
            O => \N__22120\,
            I => \N__22112\
        );

    \I__4076\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22109\
        );

    \I__4075\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22106\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__22115\,
            I => \this_ppu_M_screen_y_q_3\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__22112\,
            I => \this_ppu_M_screen_y_q_3\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__22109\,
            I => \this_ppu_M_screen_y_q_3\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__22106\,
            I => \this_ppu_M_screen_y_q_3\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22093\
        );

    \I__4069\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22090\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__22093\,
            I => \this_ppu.un3_M_screen_y_d_0_c2\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22090\,
            I => \this_ppu.un3_M_screen_y_d_0_c2\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22081\
        );

    \I__4065\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22078\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__22081\,
            I => \N__22072\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__22078\,
            I => \N__22069\
        );

    \I__4062\ : InMux
    port map (
            O => \N__22077\,
            I => \N__22066\
        );

    \I__4061\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22063\
        );

    \I__4060\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22060\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__22072\,
            I => \N__22057\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__22069\,
            I => \N__22054\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__22066\,
            I => \this_ppu_M_screen_y_q_4\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__22063\,
            I => \this_ppu_M_screen_y_q_4\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__22060\,
            I => \this_ppu_M_screen_y_q_4\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__22057\,
            I => \this_ppu_M_screen_y_q_4\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__22054\,
            I => \this_ppu_M_screen_y_q_4\
        );

    \I__4052\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22038\
        );

    \I__4051\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22035\
        );

    \I__4050\ : InMux
    port map (
            O => \N__22041\,
            I => \N__22032\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__22029\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__22035\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__22032\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__22029\,
            I => \this_ppu.M_state_qZ0Z_6\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__22022\,
            I => \this_ppu.m68_0_a2_2_cascade_\
        );

    \I__4044\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__22016\,
            I => \N__22012\
        );

    \I__4042\ : InMux
    port map (
            O => \N__22015\,
            I => \N__22009\
        );

    \I__4041\ : Span4Mux_h
    port map (
            O => \N__22012\,
            I => \N__22006\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__22009\,
            I => \N__22003\
        );

    \I__4039\ : Odrv4
    port map (
            O => \N__22006\,
            I => \this_ppu.M_state_q_ns_7\
        );

    \I__4038\ : Odrv4
    port map (
            O => \N__22003\,
            I => \this_ppu.M_state_q_ns_7\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__4036\ : InMux
    port map (
            O => \N__21995\,
            I => \N__21986\
        );

    \I__4035\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21986\
        );

    \I__4034\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21981\
        );

    \I__4033\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21981\
        );

    \I__4032\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21973\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__21986\,
            I => \N__21968\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__21981\,
            I => \N__21968\
        );

    \I__4029\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21957\
        );

    \I__4028\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21957\
        );

    \I__4027\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21957\
        );

    \I__4026\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21957\
        );

    \I__4025\ : InMux
    port map (
            O => \N__21976\,
            I => \N__21957\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__21973\,
            I => \this_ppu.N_814\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__21968\,
            I => \this_ppu.N_814\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__21957\,
            I => \this_ppu.N_814\
        );

    \I__4021\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21939\
        );

    \I__4020\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21936\
        );

    \I__4019\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21931\
        );

    \I__4018\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21931\
        );

    \I__4017\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21928\
        );

    \I__4016\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21919\
        );

    \I__4015\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21919\
        );

    \I__4014\ : InMux
    port map (
            O => \N__21943\,
            I => \N__21919\
        );

    \I__4013\ : InMux
    port map (
            O => \N__21942\,
            I => \N__21919\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__21939\,
            I => \this_ppu.N_783\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__21936\,
            I => \this_ppu.N_783\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__21931\,
            I => \this_ppu.N_783\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__21928\,
            I => \this_ppu.N_783\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__21919\,
            I => \this_ppu.N_783\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__4006\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21902\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__21902\,
            I => \this_ppu.M_state_q_RNISP3R6_3Z0Z_10\
        );

    \I__4004\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21894\
        );

    \I__4003\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21889\
        );

    \I__4002\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21889\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__21894\,
            I => \N__21886\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__21889\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__21886\,
            I => \un1_M_this_oam_address_q_c2\
        );

    \I__3998\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21878\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__3996\ : Span4Mux_h
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__21872\,
            I => \M_this_data_tmp_qZ0Z_18\
        );

    \I__3994\ : InMux
    port map (
            O => \N__21869\,
            I => \N__21866\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__21863\,
            I => \M_this_data_tmp_qZ0Z_1\
        );

    \I__3991\ : InMux
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__21854\,
            I => \M_this_data_tmp_qZ0Z_19\
        );

    \I__3988\ : CEMux
    port map (
            O => \N__21851\,
            I => \N__21845\
        );

    \I__3987\ : CEMux
    port map (
            O => \N__21850\,
            I => \N__21842\
        );

    \I__3986\ : CEMux
    port map (
            O => \N__21849\,
            I => \N__21839\
        );

    \I__3985\ : CEMux
    port map (
            O => \N__21848\,
            I => \N__21836\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21831\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__21842\,
            I => \N__21831\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21826\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__21836\,
            I => \N__21826\
        );

    \I__3980\ : Span4Mux_v
    port map (
            O => \N__21831\,
            I => \N__21821\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__21826\,
            I => \N__21818\
        );

    \I__3978\ : CEMux
    port map (
            O => \N__21825\,
            I => \N__21815\
        );

    \I__3977\ : CEMux
    port map (
            O => \N__21824\,
            I => \N__21812\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__21821\,
            I => \N_1232_0\
        );

    \I__3975\ : Odrv4
    port map (
            O => \N__21818\,
            I => \N_1232_0\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N_1232_0\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N_1232_0\
        );

    \I__3972\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__21800\,
            I => \this_ppu.M_state_q_RNISP3R6_2Z0Z_10\
        );

    \I__3970\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__21794\,
            I => \this_ppu.M_state_q_RNISP3R6_4Z0Z_10\
        );

    \I__3968\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__21788\,
            I => \this_ppu.M_state_q_RNISP3R6_0Z0Z_10\
        );

    \I__3966\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21781\
        );

    \I__3965\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21773\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__21781\,
            I => \N__21769\
        );

    \I__3963\ : InMux
    port map (
            O => \N__21780\,
            I => \N__21766\
        );

    \I__3962\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21763\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__21778\,
            I => \N__21760\
        );

    \I__3960\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21755\
        );

    \I__3959\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21755\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21752\
        );

    \I__3957\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21749\
        );

    \I__3956\ : Span4Mux_v
    port map (
            O => \N__21769\,
            I => \N__21744\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21744\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__21763\,
            I => \N__21741\
        );

    \I__3953\ : InMux
    port map (
            O => \N__21760\,
            I => \N__21738\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__21755\,
            I => \N__21735\
        );

    \I__3951\ : Odrv12
    port map (
            O => \N__21752\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__21749\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__21744\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3948\ : Odrv4
    port map (
            O => \N__21741\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__21738\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3946\ : Odrv12
    port map (
            O => \N__21735\,
            I => \this_ppu.M_state_qZ0Z_4\
        );

    \I__3945\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21718\
        );

    \I__3944\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21715\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__21718\,
            I => \N__21711\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__21715\,
            I => \N__21706\
        );

    \I__3941\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21703\
        );

    \I__3940\ : Span4Mux_v
    port map (
            O => \N__21711\,
            I => \N__21700\
        );

    \I__3939\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21695\
        );

    \I__3938\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21695\
        );

    \I__3937\ : Span4Mux_h
    port map (
            O => \N__21706\,
            I => \N__21690\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21690\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__21700\,
            I => \N__21685\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__21695\,
            I => \N__21685\
        );

    \I__3933\ : Sp12to4
    port map (
            O => \N__21690\,
            I => \N__21682\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__21685\,
            I => \N__21679\
        );

    \I__3931\ : Odrv12
    port map (
            O => \N__21682\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__21679\,
            I => \this_ppu.M_state_qZ0Z_10\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__21674\,
            I => \this_ppu.N_835_0_cascade_\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__21671\,
            I => \this_ppu.N_783_cascade_\
        );

    \I__3927\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__21665\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__3923\ : Span4Mux_v
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__21650\,
            I => \this_ppu.oam_cache.mem_2\
        );

    \I__3920\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21640\
        );

    \I__3918\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21636\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__21640\,
            I => \N__21633\
        );

    \I__3916\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21630\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__21636\,
            I => \this_ppu.N_60_0\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__21633\,
            I => \this_ppu.N_60_0\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__21630\,
            I => \this_ppu.N_60_0\
        );

    \I__3912\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21617\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__21622\,
            I => \N__21614\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__21621\,
            I => \N__21609\
        );

    \I__3909\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21605\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21602\
        );

    \I__3907\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21595\
        );

    \I__3906\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21595\
        );

    \I__3905\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21595\
        );

    \I__3904\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21591\
        );

    \I__3903\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21588\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__21605\,
            I => \N__21585\
        );

    \I__3901\ : Span4Mux_v
    port map (
            O => \N__21602\,
            I => \N__21580\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__21595\,
            I => \N__21580\
        );

    \I__3899\ : InMux
    port map (
            O => \N__21594\,
            I => \N__21576\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__21591\,
            I => \N__21571\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21571\
        );

    \I__3896\ : Span4Mux_h
    port map (
            O => \N__21585\,
            I => \N__21562\
        );

    \I__3895\ : Span4Mux_h
    port map (
            O => \N__21580\,
            I => \N__21562\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21559\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__21576\,
            I => \N__21554\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__21571\,
            I => \N__21554\
        );

    \I__3891\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21551\
        );

    \I__3890\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21548\
        );

    \I__3889\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21543\
        );

    \I__3888\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21543\
        );

    \I__3887\ : Sp12to4
    port map (
            O => \N__21562\,
            I => \N__21538\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__21559\,
            I => \N__21538\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__21554\,
            I => \N__21535\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__21551\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__21548\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__21543\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__21538\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__21535\,
            I => \this_ppu.M_state_qZ0Z_0\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__21524\,
            I => \N__21516\
        );

    \I__3878\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21507\
        );

    \I__3877\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21507\
        );

    \I__3876\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21507\
        );

    \I__3875\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21507\
        );

    \I__3874\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21501\
        );

    \I__3873\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21498\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__21507\,
            I => \N__21495\
        );

    \I__3871\ : InMux
    port map (
            O => \N__21506\,
            I => \N__21492\
        );

    \I__3870\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21489\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21486\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__21501\,
            I => \N__21483\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__21498\,
            I => \N__21480\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__21495\,
            I => \N__21477\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__21492\,
            I => \N__21473\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__21489\,
            I => \N__21468\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__21486\,
            I => \N__21468\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__21483\,
            I => \N__21465\
        );

    \I__3861\ : Span4Mux_h
    port map (
            O => \N__21480\,
            I => \N__21460\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__21477\,
            I => \N__21460\
        );

    \I__3859\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21457\
        );

    \I__3858\ : Span4Mux_h
    port map (
            O => \N__21473\,
            I => \N__21454\
        );

    \I__3857\ : Span4Mux_h
    port map (
            O => \N__21468\,
            I => \N__21449\
        );

    \I__3856\ : Span4Mux_v
    port map (
            O => \N__21465\,
            I => \N__21449\
        );

    \I__3855\ : Odrv4
    port map (
            O => \N__21460\,
            I => \this_ppu.N_835_0\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__21457\,
            I => \this_ppu.N_835_0\
        );

    \I__3853\ : Odrv4
    port map (
            O => \N__21454\,
            I => \this_ppu.N_835_0\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__21449\,
            I => \this_ppu.N_835_0\
        );

    \I__3851\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21431\
        );

    \I__3850\ : InMux
    port map (
            O => \N__21439\,
            I => \N__21428\
        );

    \I__3849\ : InMux
    port map (
            O => \N__21438\,
            I => \N__21417\
        );

    \I__3848\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21417\
        );

    \I__3847\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21417\
        );

    \I__3846\ : InMux
    port map (
            O => \N__21435\,
            I => \N__21417\
        );

    \I__3845\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21417\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__21431\,
            I => \N__21414\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__21428\,
            I => \N__21409\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21409\
        );

    \I__3841\ : Span4Mux_v
    port map (
            O => \N__21414\,
            I => \N__21406\
        );

    \I__3840\ : Span4Mux_h
    port map (
            O => \N__21409\,
            I => \N__21403\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__21406\,
            I => \this_ppu.N_807\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__21403\,
            I => \this_ppu.N_807\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__21398\,
            I => \N__21395\
        );

    \I__3836\ : InMux
    port map (
            O => \N__21395\,
            I => \N__21392\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21389\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__21389\,
            I => \N__21386\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__21386\,
            I => \M_this_scroll_qZ0Z_8\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__21383\,
            I => \N_829_0_cascade_\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__21380\,
            I => \N_58_0_cascade_\
        );

    \I__3830\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21369\
        );

    \I__3829\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21366\
        );

    \I__3828\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21363\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \N__21360\
        );

    \I__3826\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21356\
        );

    \I__3825\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21353\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__21369\,
            I => \N__21350\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__21366\,
            I => \N__21345\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__21363\,
            I => \N__21345\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21342\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__21359\,
            I => \N__21338\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21335\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__21353\,
            I => \N__21332\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__21350\,
            I => \N__21327\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__21345\,
            I => \N__21327\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__21342\,
            I => \N__21324\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21321\
        );

    \I__3813\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21318\
        );

    \I__3812\ : Odrv4
    port map (
            O => \N__21335\,
            I => \this_ppu.N_97_mux\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__21332\,
            I => \this_ppu.N_97_mux\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__21327\,
            I => \this_ppu.N_97_mux\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__21324\,
            I => \this_ppu.N_97_mux\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__21321\,
            I => \this_ppu.N_97_mux\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__21318\,
            I => \this_ppu.N_97_mux\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__21305\,
            I => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_\
        );

    \I__3805\ : InMux
    port map (
            O => \N__21302\,
            I => \N__21299\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__21299\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__21296\,
            I => \N__21292\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21289\
        );

    \I__3801\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21286\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__21286\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_2\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__21283\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_2\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__3796\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21271\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21268\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__21271\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_1\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__21268\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_1\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__21263\,
            I => \N__21259\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__21262\,
            I => \N__21256\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21253\
        );

    \I__3789\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21250\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21247\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__21250\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_7\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__21247\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_7\
        );

    \I__3785\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__21239\,
            I => \this_ppu.m9_0_a2_4\
        );

    \I__3783\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21232\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__21235\,
            I => \N__21228\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21225\
        );

    \I__3780\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21222\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21228\,
            I => \N__21219\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__21225\,
            I => \N__21214\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21214\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__21219\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_0\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__21214\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_0\
        );

    \I__3774\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__21206\,
            I => \N__21203\
        );

    \I__3772\ : Span4Mux_v
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__21200\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_axb_0\
        );

    \I__3770\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__21194\,
            I => \this_ppu.un1_M_surface_x_q_c2\
        );

    \I__3768\ : InMux
    port map (
            O => \N__21191\,
            I => \N__21183\
        );

    \I__3767\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21183\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21189\,
            I => \N__21180\
        );

    \I__3765\ : InMux
    port map (
            O => \N__21188\,
            I => \N__21177\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21183\,
            I => \this_ppu.M_oam_curr_dZ0Z25\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__21180\,
            I => \this_ppu.M_oam_curr_dZ0Z25\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__21177\,
            I => \this_ppu.M_oam_curr_dZ0Z25\
        );

    \I__3761\ : InMux
    port map (
            O => \N__21170\,
            I => \N__21167\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__21167\,
            I => \N__21160\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__21166\,
            I => \N__21157\
        );

    \I__3758\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21152\
        );

    \I__3757\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21149\
        );

    \I__3756\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21146\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__21160\,
            I => \N__21143\
        );

    \I__3754\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21140\
        );

    \I__3753\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21135\
        );

    \I__3752\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21135\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__21130\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__21149\,
            I => \N__21130\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__21146\,
            I => \N__21127\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__21143\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__21140\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__21135\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__21130\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__21127\,
            I => \this_ppu.M_state_qZ0Z_7\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__21116\,
            I => \N__21109\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__21115\,
            I => \N__21106\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21103\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21100\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21092\
        );

    \I__3738\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21092\
        );

    \I__3737\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21092\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__21103\,
            I => \N__21086\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21086\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21083\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21080\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21077\
        );

    \I__3731\ : Span4Mux_v
    port map (
            O => \N__21086\,
            I => \N__21074\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__21083\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__3729\ : Odrv4
    port map (
            O => \N__21080\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__21077\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__3727\ : Odrv4
    port map (
            O => \N__21074\,
            I => \this_ppu.M_state_qZ0Z_9\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__21065\,
            I => \this_ppu.un1_M_surface_x_q_c1_cascade_\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__21062\,
            I => \N__21059\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__21053\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__21053\,
            I => \M_this_scroll_qZ0Z_10\
        );

    \I__3721\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__21044\,
            I => \M_this_scroll_qZ0Z_11\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__21038\,
            I => \M_this_scroll_qZ0Z_13\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21032\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__3714\ : Span4Mux_v
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__3713\ : Odrv4
    port map (
            O => \N__21026\,
            I => \M_this_scroll_qZ0Z_14\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__21023\,
            I => \this_ppu.N_798_0_cascade_\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__21020\,
            I => \N__21017\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__21014\,
            I => \this_ppu.un1_M_surface_x_q_c3\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__21011\,
            I => \this_ppu.un1_M_surface_x_q_c3_cascade_\
        );

    \I__3707\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__21005\,
            I => \this_ppu.N_798_0\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__21002\,
            I => \this_ppu.un1_M_surface_x_q_c2_cascade_\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__20999\,
            I => \this_ppu.un1_M_surface_x_q_c5_cascade_\
        );

    \I__3703\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20989\
        );

    \I__3701\ : InMux
    port map (
            O => \N__20992\,
            I => \N__20986\
        );

    \I__3700\ : Odrv4
    port map (
            O => \N__20989\,
            I => \this_ppu.N_800\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__20986\,
            I => \this_ppu.N_800\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__20981\,
            I => \this_ppu.N_800_cascade_\
        );

    \I__3697\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20972\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__20977\,
            I => \N__20968\
        );

    \I__3695\ : InMux
    port map (
            O => \N__20976\,
            I => \N__20965\
        );

    \I__3694\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20962\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__20972\,
            I => \N__20959\
        );

    \I__3692\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20956\
        );

    \I__3691\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20953\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20948\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__20962\,
            I => \N__20948\
        );

    \I__3688\ : Span4Mux_v
    port map (
            O => \N__20959\,
            I => \N__20941\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20941\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__20953\,
            I => \N__20941\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__20948\,
            I => \N__20938\
        );

    \I__3684\ : Span4Mux_v
    port map (
            O => \N__20941\,
            I => \N__20935\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__20938\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__20935\,
            I => \this_ppu.M_state_qZ0Z_11\
        );

    \I__3681\ : CEMux
    port map (
            O => \N__20930\,
            I => \N__20927\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20924\
        );

    \I__3679\ : Span4Mux_v
    port map (
            O => \N__20924\,
            I => \N__20921\
        );

    \I__3678\ : Span4Mux_h
    port map (
            O => \N__20921\,
            I => \N__20918\
        );

    \I__3677\ : Odrv4
    port map (
            O => \N__20918\,
            I => \N_18\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__20915\,
            I => \this_ppu.un3_M_screen_y_d_0_c4_cascade_\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__20912\,
            I => \N__20909\
        );

    \I__3674\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__20900\,
            I => \this_ppu.N_802\
        );

    \I__3670\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20894\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__3668\ : Span12Mux_h
    port map (
            O => \N__20891\,
            I => \N__20888\
        );

    \I__3667\ : Span12Mux_v
    port map (
            O => \N__20888\,
            I => \N__20885\
        );

    \I__3666\ : Odrv12
    port map (
            O => \N__20885\,
            I => \this_spr_ram.mem_out_bus7_3\
        );

    \I__3665\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__3663\ : Span12Mux_v
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__3662\ : Span12Mux_h
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__3661\ : Odrv12
    port map (
            O => \N__20870\,
            I => \this_spr_ram.mem_out_bus3_3\
        );

    \I__3660\ : InMux
    port map (
            O => \N__20867\,
            I => \N__20860\
        );

    \I__3659\ : InMux
    port map (
            O => \N__20866\,
            I => \N__20853\
        );

    \I__3658\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20853\
        );

    \I__3657\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20853\
        );

    \I__3656\ : InMux
    port map (
            O => \N__20863\,
            I => \N__20849\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__20860\,
            I => \N__20844\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20844\
        );

    \I__3653\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20841\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__20849\,
            I => \N__20831\
        );

    \I__3651\ : Span4Mux_v
    port map (
            O => \N__20844\,
            I => \N__20831\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__20841\,
            I => \N__20831\
        );

    \I__3649\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20819\
        );

    \I__3648\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20819\
        );

    \I__3647\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20816\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__20831\,
            I => \N__20813\
        );

    \I__3645\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20806\
        );

    \I__3644\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20806\
        );

    \I__3643\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20806\
        );

    \I__3642\ : InMux
    port map (
            O => \N__20827\,
            I => \N__20801\
        );

    \I__3641\ : InMux
    port map (
            O => \N__20826\,
            I => \N__20801\
        );

    \I__3640\ : InMux
    port map (
            O => \N__20825\,
            I => \N__20798\
        );

    \I__3639\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20795\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__20819\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__20816\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__20813\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__20806\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__20801\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__20798\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__20795\,
            I => \this_spr_ram.mem_radregZ0Z_13\
        );

    \I__3631\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__3629\ : Odrv4
    port map (
            O => \N__20774\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\
        );

    \I__3628\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20764\
        );

    \I__3627\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20761\
        );

    \I__3626\ : InMux
    port map (
            O => \N__20769\,
            I => \N__20756\
        );

    \I__3625\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20756\
        );

    \I__3624\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20753\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20750\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__20761\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__20756\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__20753\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__3619\ : Odrv12
    port map (
            O => \N__20750\,
            I => \this_ppu.M_state_qZ0Z_5\
        );

    \I__3618\ : CascadeMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__3617\ : InMux
    port map (
            O => \N__20738\,
            I => \N__20734\
        );

    \I__3616\ : InMux
    port map (
            O => \N__20737\,
            I => \N__20731\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__20734\,
            I => \N__20726\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20726\
        );

    \I__3613\ : Span4Mux_v
    port map (
            O => \N__20726\,
            I => \N__20723\
        );

    \I__3612\ : Span4Mux_h
    port map (
            O => \N__20723\,
            I => \N__20720\
        );

    \I__3611\ : Span4Mux_v
    port map (
            O => \N__20720\,
            I => \N__20717\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__20717\,
            I => \this_ppu.N_796_0\
        );

    \I__3609\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__20711\,
            I => \this_ppu.M_state_qZ0Z_8\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__20708\,
            I => \this_ppu.un1_M_surface_x_q_c6_cascade_\
        );

    \I__3606\ : InMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__20702\,
            I => \N__20699\
        );

    \I__3604\ : Span12Mux_v
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__3603\ : Span12Mux_h
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__3602\ : Odrv12
    port map (
            O => \N__20693\,
            I => \M_this_map_ram_read_data_7\
        );

    \I__3601\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__20687\,
            I => \N__20684\
        );

    \I__3599\ : Odrv12
    port map (
            O => \N__20684\,
            I => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20678\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__20678\,
            I => \N__20675\
        );

    \I__3596\ : Span4Mux_h
    port map (
            O => \N__20675\,
            I => \N__20672\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__20672\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_3\
        );

    \I__3594\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20666\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20663\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__3591\ : Span4Mux_h
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__3590\ : Sp12to4
    port map (
            O => \N__20657\,
            I => \N__20654\
        );

    \I__3589\ : Span12Mux_v
    port map (
            O => \N__20654\,
            I => \N__20651\
        );

    \I__3588\ : Odrv12
    port map (
            O => \N__20651\,
            I => \M_this_map_ram_read_data_3\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__20648\,
            I => \N__20644\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__20647\,
            I => \N__20641\
        );

    \I__3585\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20634\
        );

    \I__3584\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20631\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__20640\,
            I => \N__20628\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__20639\,
            I => \N__20624\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__20638\,
            I => \N__20616\
        );

    \I__3580\ : CascadeMux
    port map (
            O => \N__20637\,
            I => \N__20613\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20607\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__20631\,
            I => \N__20607\
        );

    \I__3577\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20604\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__20627\,
            I => \N__20601\
        );

    \I__3575\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20598\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__20623\,
            I => \N__20595\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__20622\,
            I => \N__20592\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__20621\,
            I => \N__20589\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__20620\,
            I => \N__20585\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__20619\,
            I => \N__20582\
        );

    \I__3569\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20577\
        );

    \I__3568\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20574\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__20612\,
            I => \N__20571\
        );

    \I__3566\ : Span4Mux_s2_v
    port map (
            O => \N__20607\,
            I => \N__20566\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20566\
        );

    \I__3564\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20563\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20560\
        );

    \I__3562\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20557\
        );

    \I__3561\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20554\
        );

    \I__3560\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20551\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__20588\,
            I => \N__20548\
        );

    \I__3558\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20545\
        );

    \I__3557\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20542\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__20581\,
            I => \N__20539\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__20580\,
            I => \N__20536\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20533\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20530\
        );

    \I__3552\ : InMux
    port map (
            O => \N__20571\,
            I => \N__20527\
        );

    \I__3551\ : Span4Mux_v
    port map (
            O => \N__20566\,
            I => \N__20522\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20522\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__20560\,
            I => \N__20517\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20517\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__20554\,
            I => \N__20514\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20511\
        );

    \I__3545\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20508\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__20545\,
            I => \N__20503\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20503\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20500\
        );

    \I__3541\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20497\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__20533\,
            I => \N__20492\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__20530\,
            I => \N__20492\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__20527\,
            I => \N__20489\
        );

    \I__3537\ : Span4Mux_h
    port map (
            O => \N__20522\,
            I => \N__20486\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__20517\,
            I => \N__20477\
        );

    \I__3535\ : Span4Mux_v
    port map (
            O => \N__20514\,
            I => \N__20477\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__20511\,
            I => \N__20477\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20477\
        );

    \I__3532\ : Span4Mux_s2_v
    port map (
            O => \N__20503\,
            I => \N__20472\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__20500\,
            I => \N__20472\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__20497\,
            I => \N__20469\
        );

    \I__3529\ : Sp12to4
    port map (
            O => \N__20492\,
            I => \N__20464\
        );

    \I__3528\ : Span12Mux_s8_h
    port map (
            O => \N__20489\,
            I => \N__20464\
        );

    \I__3527\ : Span4Mux_v
    port map (
            O => \N__20486\,
            I => \N__20459\
        );

    \I__3526\ : Span4Mux_h
    port map (
            O => \N__20477\,
            I => \N__20459\
        );

    \I__3525\ : Span4Mux_v
    port map (
            O => \N__20472\,
            I => \N__20454\
        );

    \I__3524\ : Span4Mux_h
    port map (
            O => \N__20469\,
            I => \N__20454\
        );

    \I__3523\ : Span12Mux_v
    port map (
            O => \N__20464\,
            I => \N__20449\
        );

    \I__3522\ : Sp12to4
    port map (
            O => \N__20459\,
            I => \N__20449\
        );

    \I__3521\ : Span4Mux_h
    port map (
            O => \N__20454\,
            I => \N__20446\
        );

    \I__3520\ : Odrv12
    port map (
            O => \N__20449\,
            I => \M_this_ppu_spr_addr_9\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__20446\,
            I => \M_this_ppu_spr_addr_9\
        );

    \I__3518\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__3516\ : Span4Mux_h
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__3515\ : Odrv4
    port map (
            O => \N__20432\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_4\
        );

    \I__3514\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20426\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20423\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__20423\,
            I => \N__20420\
        );

    \I__3511\ : Span4Mux_v
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__3510\ : Sp12to4
    port map (
            O => \N__20417\,
            I => \N__20414\
        );

    \I__3509\ : Span12Mux_h
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__3508\ : Span12Mux_v
    port map (
            O => \N__20411\,
            I => \N__20408\
        );

    \I__3507\ : Odrv12
    port map (
            O => \N__20408\,
            I => \M_this_map_ram_read_data_4\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__20405\,
            I => \N__20402\
        );

    \I__3505\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20397\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__20401\,
            I => \N__20394\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__20400\,
            I => \N__20390\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__20397\,
            I => \N__20386\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20383\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__20393\,
            I => \N__20380\
        );

    \I__3499\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20374\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__20389\,
            I => \N__20371\
        );

    \I__3497\ : Span4Mux_s2_v
    port map (
            O => \N__20386\,
            I => \N__20366\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__20383\,
            I => \N__20366\
        );

    \I__3495\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20363\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__20379\,
            I => \N__20360\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__20378\,
            I => \N__20356\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__20377\,
            I => \N__20353\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20347\
        );

    \I__3490\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20344\
        );

    \I__3489\ : Span4Mux_h
    port map (
            O => \N__20366\,
            I => \N__20338\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__20363\,
            I => \N__20338\
        );

    \I__3487\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20335\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__20359\,
            I => \N__20332\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20329\
        );

    \I__3484\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20326\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__20352\,
            I => \N__20323\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__20351\,
            I => \N__20319\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__20350\,
            I => \N__20316\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__20347\,
            I => \N__20309\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__20344\,
            I => \N__20309\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__20343\,
            I => \N__20306\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__20338\,
            I => \N__20301\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20301\
        );

    \I__3475\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20298\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__20329\,
            I => \N__20295\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20292\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20289\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__20322\,
            I => \N__20286\
        );

    \I__3470\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20283\
        );

    \I__3469\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20280\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__20315\,
            I => \N__20277\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__20314\,
            I => \N__20274\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__20309\,
            I => \N__20271\
        );

    \I__3465\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20268\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__20301\,
            I => \N__20263\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20263\
        );

    \I__3462\ : Span4Mux_v
    port map (
            O => \N__20295\,
            I => \N__20256\
        );

    \I__3461\ : Span4Mux_h
    port map (
            O => \N__20292\,
            I => \N__20256\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20256\
        );

    \I__3459\ : InMux
    port map (
            O => \N__20286\,
            I => \N__20253\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__20283\,
            I => \N__20248\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__20280\,
            I => \N__20248\
        );

    \I__3456\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20245\
        );

    \I__3455\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20242\
        );

    \I__3454\ : Sp12to4
    port map (
            O => \N__20271\,
            I => \N__20237\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__20268\,
            I => \N__20237\
        );

    \I__3452\ : Span4Mux_v
    port map (
            O => \N__20263\,
            I => \N__20230\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__20256\,
            I => \N__20230\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__20253\,
            I => \N__20230\
        );

    \I__3449\ : Span4Mux_s2_v
    port map (
            O => \N__20248\,
            I => \N__20225\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__20245\,
            I => \N__20225\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20222\
        );

    \I__3446\ : Span12Mux_h
    port map (
            O => \N__20237\,
            I => \N__20219\
        );

    \I__3445\ : Sp12to4
    port map (
            O => \N__20230\,
            I => \N__20216\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__20225\,
            I => \N__20211\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__20222\,
            I => \N__20211\
        );

    \I__3442\ : Span12Mux_v
    port map (
            O => \N__20219\,
            I => \N__20206\
        );

    \I__3441\ : Span12Mux_h
    port map (
            O => \N__20216\,
            I => \N__20206\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__20211\,
            I => \N__20203\
        );

    \I__3439\ : Odrv12
    port map (
            O => \N__20206\,
            I => \M_this_ppu_spr_addr_10\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__20203\,
            I => \M_this_ppu_spr_addr_10\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__20198\,
            I => \N__20193\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__20197\,
            I => \N__20189\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__20196\,
            I => \N__20186\
        );

    \I__3434\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20182\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__20192\,
            I => \N__20179\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20173\
        );

    \I__3431\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20170\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__20185\,
            I => \N__20166\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20162\
        );

    \I__3428\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20159\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__20178\,
            I => \N__20156\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__20177\,
            I => \N__20152\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__20176\,
            I => \N__20149\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__20173\,
            I => \N__20140\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__20170\,
            I => \N__20140\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__20169\,
            I => \N__20137\
        );

    \I__3421\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20134\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__20165\,
            I => \N__20131\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__20162\,
            I => \N__20126\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__20159\,
            I => \N__20126\
        );

    \I__3417\ : InMux
    port map (
            O => \N__20156\,
            I => \N__20123\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__20155\,
            I => \N__20120\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20116\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20113\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__20148\,
            I => \N__20110\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__20147\,
            I => \N__20107\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__20146\,
            I => \N__20104\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__20145\,
            I => \N__20101\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__20140\,
            I => \N__20098\
        );

    \I__3408\ : InMux
    port map (
            O => \N__20137\,
            I => \N__20095\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__20134\,
            I => \N__20092\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20089\
        );

    \I__3405\ : Span4Mux_h
    port map (
            O => \N__20126\,
            I => \N__20084\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20084\
        );

    \I__3403\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20081\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__20119\,
            I => \N__20078\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__20116\,
            I => \N__20073\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20073\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20070\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20067\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20104\,
            I => \N__20064\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20061\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__20098\,
            I => \N__20058\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20095\,
            I => \N__20055\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__20092\,
            I => \N__20046\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__20089\,
            I => \N__20046\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__20084\,
            I => \N__20046\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20046\
        );

    \I__3389\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20043\
        );

    \I__3388\ : Span4Mux_s2_v
    port map (
            O => \N__20073\,
            I => \N__20038\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__20070\,
            I => \N__20038\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20035\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20030\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__20061\,
            I => \N__20030\
        );

    \I__3383\ : Sp12to4
    port map (
            O => \N__20058\,
            I => \N__20025\
        );

    \I__3382\ : Span12Mux_h
    port map (
            O => \N__20055\,
            I => \N__20025\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__20046\,
            I => \N__20022\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__20019\
        );

    \I__3379\ : Span4Mux_v
    port map (
            O => \N__20038\,
            I => \N__20014\
        );

    \I__3378\ : Span4Mux_h
    port map (
            O => \N__20035\,
            I => \N__20014\
        );

    \I__3377\ : Span12Mux_s10_v
    port map (
            O => \N__20030\,
            I => \N__20005\
        );

    \I__3376\ : Span12Mux_v
    port map (
            O => \N__20025\,
            I => \N__20005\
        );

    \I__3375\ : Sp12to4
    port map (
            O => \N__20022\,
            I => \N__20005\
        );

    \I__3374\ : Span12Mux_s7_h
    port map (
            O => \N__20019\,
            I => \N__20005\
        );

    \I__3373\ : Span4Mux_h
    port map (
            O => \N__20014\,
            I => \N__20002\
        );

    \I__3372\ : Odrv12
    port map (
            O => \N__20005\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__20002\,
            I => \M_this_ppu_spr_addr_0\
        );

    \I__3370\ : InMux
    port map (
            O => \N__19997\,
            I => \N__19994\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__19994\,
            I => \N__19991\
        );

    \I__3368\ : Span12Mux_h
    port map (
            O => \N__19991\,
            I => \N__19988\
        );

    \I__3367\ : Span12Mux_v
    port map (
            O => \N__19988\,
            I => \N__19985\
        );

    \I__3366\ : Odrv12
    port map (
            O => \N__19985\,
            I => \this_spr_ram.mem_out_bus6_3\
        );

    \I__3365\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19979\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__19979\,
            I => \N__19976\
        );

    \I__3363\ : Span12Mux_v
    port map (
            O => \N__19976\,
            I => \N__19973\
        );

    \I__3362\ : Span12Mux_h
    port map (
            O => \N__19973\,
            I => \N__19970\
        );

    \I__3361\ : Odrv12
    port map (
            O => \N__19970\,
            I => \this_spr_ram.mem_out_bus2_3\
        );

    \I__3360\ : InMux
    port map (
            O => \N__19967\,
            I => \N__19964\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__19964\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\
        );

    \I__3358\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__19958\,
            I => \N__19955\
        );

    \I__3356\ : Span4Mux_h
    port map (
            O => \N__19955\,
            I => \N__19952\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__19952\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_5\
        );

    \I__3354\ : InMux
    port map (
            O => \N__19949\,
            I => \N__19946\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__19946\,
            I => \N__19943\
        );

    \I__3352\ : Span4Mux_h
    port map (
            O => \N__19943\,
            I => \N__19940\
        );

    \I__3351\ : Sp12to4
    port map (
            O => \N__19940\,
            I => \N__19937\
        );

    \I__3350\ : Span12Mux_v
    port map (
            O => \N__19937\,
            I => \N__19934\
        );

    \I__3349\ : Span12Mux_h
    port map (
            O => \N__19934\,
            I => \N__19931\
        );

    \I__3348\ : Odrv12
    port map (
            O => \N__19931\,
            I => \M_this_map_ram_read_data_5\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__19928\,
            I => \N__19922\
        );

    \I__3346\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19919\
        );

    \I__3345\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19916\
        );

    \I__3344\ : InMux
    port map (
            O => \N__19925\,
            I => \N__19912\
        );

    \I__3343\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19907\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19903\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19900\
        );

    \I__3340\ : InMux
    port map (
            O => \N__19915\,
            I => \N__19897\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19894\
        );

    \I__3338\ : InMux
    port map (
            O => \N__19911\,
            I => \N__19891\
        );

    \I__3337\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19888\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__19907\,
            I => \N__19885\
        );

    \I__3335\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19882\
        );

    \I__3334\ : Span4Mux_h
    port map (
            O => \N__19903\,
            I => \N__19875\
        );

    \I__3333\ : Span4Mux_v
    port map (
            O => \N__19900\,
            I => \N__19875\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__19897\,
            I => \N__19875\
        );

    \I__3331\ : Span4Mux_h
    port map (
            O => \N__19894\,
            I => \N__19872\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19869\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__19888\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3328\ : Odrv12
    port map (
            O => \N__19885\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__19882\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__19875\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__19872\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__19869\,
            I => \this_spr_ram.mem_radregZ0Z_11\
        );

    \I__3323\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__19853\,
            I => \this_ppu.N_797\
        );

    \I__3321\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__19847\,
            I => \M_this_data_tmp_qZ0Z_2\
        );

    \I__3319\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19841\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__19838\,
            I => \M_this_data_tmp_qZ0Z_21\
        );

    \I__3316\ : InMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__19832\,
            I => \N__19829\
        );

    \I__3314\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19826\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__19826\,
            I => \N__19823\
        );

    \I__3312\ : Span4Mux_v
    port map (
            O => \N__19823\,
            I => \N__19820\
        );

    \I__3311\ : Span4Mux_v
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__19817\,
            I => \N__19814\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__19814\,
            I => \this_spr_ram.mem_out_bus7_0\
        );

    \I__3308\ : InMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19805\
        );

    \I__3306\ : Span4Mux_h
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__19796\,
            I => \this_spr_ram.mem_out_bus3_0\
        );

    \I__3302\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__3300\ : Span12Mux_v
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3299\ : Span12Mux_h
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__3298\ : Odrv12
    port map (
            O => \N__19781\,
            I => \this_spr_ram.mem_out_bus4_0\
        );

    \I__3297\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__3295\ : Span4Mux_v
    port map (
            O => \N__19772\,
            I => \N__19769\
        );

    \I__3294\ : Span4Mux_h
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__19766\,
            I => \this_spr_ram.mem_out_bus0_0\
        );

    \I__3292\ : InMux
    port map (
            O => \N__19763\,
            I => \N__19760\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19757\
        );

    \I__3290\ : Span4Mux_h
    port map (
            O => \N__19757\,
            I => \N__19754\
        );

    \I__3289\ : Span4Mux_v
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__3288\ : Span4Mux_h
    port map (
            O => \N__19751\,
            I => \N__19748\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__19745\,
            I => \this_spr_ram.mem_out_bus5_0\
        );

    \I__3285\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19739\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__19730\,
            I => \this_spr_ram.mem_out_bus1_0\
        );

    \I__3280\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19724\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__3278\ : Sp12to4
    port map (
            O => \N__19721\,
            I => \N__19718\
        );

    \I__3277\ : Span12Mux_v
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__3276\ : Span12Mux_h
    port map (
            O => \N__19715\,
            I => \N__19712\
        );

    \I__3275\ : Odrv12
    port map (
            O => \N__19712\,
            I => \this_spr_ram.mem_out_bus6_0\
        );

    \I__3274\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19706\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19703\
        );

    \I__3272\ : Span12Mux_v
    port map (
            O => \N__19703\,
            I => \N__19700\
        );

    \I__3271\ : Span12Mux_h
    port map (
            O => \N__19700\,
            I => \N__19697\
        );

    \I__3270\ : Odrv12
    port map (
            O => \N__19697\,
            I => \this_spr_ram.mem_out_bus2_0\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__19694\,
            I => \N__19689\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__19693\,
            I => \N__19686\
        );

    \I__3267\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19683\
        );

    \I__3266\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19679\
        );

    \I__3265\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19676\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__19683\,
            I => \N__19673\
        );

    \I__3263\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19670\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19665\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19665\
        );

    \I__3260\ : Span4Mux_v
    port map (
            O => \N__19673\,
            I => \N__19662\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__19670\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__3258\ : Odrv12
    port map (
            O => \N__19665\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__3257\ : Odrv4
    port map (
            O => \N__19662\,
            I => \this_spr_ram.mem_radregZ0Z_12\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__19655\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\
        );

    \I__3255\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__19649\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\
        );

    \I__3253\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__19643\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\
        );

    \I__3251\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__19637\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\
        );

    \I__3249\ : InMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__19631\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19624\
        );

    \I__3246\ : InMux
    port map (
            O => \N__19627\,
            I => \N__19621\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__3243\ : Span4Mux_v
    port map (
            O => \N__19618\,
            I => \N__19612\
        );

    \I__3242\ : Span4Mux_v
    port map (
            O => \N__19615\,
            I => \N__19609\
        );

    \I__3241\ : Odrv4
    port map (
            O => \N__19612\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__3240\ : Odrv4
    port map (
            O => \N__19609\,
            I => \M_this_spr_ram_read_data_0\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__19604\,
            I => \N__19601\
        );

    \I__3238\ : CascadeBuf
    port map (
            O => \N__19601\,
            I => \N__19598\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__19598\,
            I => \N__19595\
        );

    \I__3236\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19591\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__19594\,
            I => \N__19588\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__19591\,
            I => \N__19584\
        );

    \I__3233\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19581\
        );

    \I__3232\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19578\
        );

    \I__3231\ : Span12Mux_s7_v
    port map (
            O => \N__19584\,
            I => \N__19575\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__19581\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__19578\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__3228\ : Odrv12
    port map (
            O => \N__19575\,
            I => \M_this_oam_address_qZ0Z_3\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__3226\ : CascadeBuf
    port map (
            O => \N__19565\,
            I => \N__19562\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__19562\,
            I => \N__19559\
        );

    \I__3224\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19556\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__19553\,
            I => \N__19547\
        );

    \I__3221\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19542\
        );

    \I__3220\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19542\
        );

    \I__3219\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19539\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__19547\,
            I => \N__19536\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__19542\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__19539\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__3215\ : Odrv4
    port map (
            O => \N__19536\,
            I => \M_this_oam_address_qZ0Z_2\
        );

    \I__3214\ : InMux
    port map (
            O => \N__19529\,
            I => \N__19523\
        );

    \I__3213\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19523\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__19523\,
            I => \un1_M_this_oam_address_q_c4\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__19520\,
            I => \N__19517\
        );

    \I__3210\ : CascadeBuf
    port map (
            O => \N__19517\,
            I => \N__19514\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__3208\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19505\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__19505\,
            I => \N__19500\
        );

    \I__3205\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19497\
        );

    \I__3204\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19494\
        );

    \I__3203\ : Span4Mux_v
    port map (
            O => \N__19500\,
            I => \N__19491\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__19497\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__19494\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__19491\,
            I => \M_this_oam_address_qZ0Z_5\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \un1_M_this_oam_address_q_c4_cascade_\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__3197\ : CascadeBuf
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \N__19472\
        );

    \I__3195\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19469\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__19469\,
            I => \N__19465\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__3192\ : Span4Mux_h
    port map (
            O => \N__19465\,
            I => \N__19457\
        );

    \I__3191\ : InMux
    port map (
            O => \N__19462\,
            I => \N__19454\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19461\,
            I => \N__19451\
        );

    \I__3189\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19448\
        );

    \I__3188\ : Span4Mux_v
    port map (
            O => \N__19457\,
            I => \N__19445\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__19454\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__19451\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__19448\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__19445\,
            I => \M_this_oam_address_qZ0Z_4\
        );

    \I__3183\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19430\
        );

    \I__3182\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19430\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__19430\,
            I => \un1_M_this_oam_address_q_c6\
        );

    \I__3180\ : CEMux
    port map (
            O => \N__19427\,
            I => \N__19423\
        );

    \I__3179\ : CEMux
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__19417\,
            I => \N_1240_0\
        );

    \I__3175\ : Odrv12
    port map (
            O => \N__19414\,
            I => \N_1240_0\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__19409\,
            I => \M_this_oam_ram_write_data_0_sqmuxa_cascade_\
        );

    \I__3173\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19403\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19400\
        );

    \I__3171\ : Span4Mux_s2_v
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__3170\ : Span4Mux_h
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__19394\,
            I => \M_this_oam_ram_write_data_26\
        );

    \I__3168\ : CEMux
    port map (
            O => \N__19391\,
            I => \N__19387\
        );

    \I__3167\ : CEMux
    port map (
            O => \N__19390\,
            I => \N__19366\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__19387\,
            I => \N__19359\
        );

    \I__3165\ : InMux
    port map (
            O => \N__19386\,
            I => \N__19352\
        );

    \I__3164\ : InMux
    port map (
            O => \N__19385\,
            I => \N__19352\
        );

    \I__3163\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19352\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19341\
        );

    \I__3161\ : InMux
    port map (
            O => \N__19382\,
            I => \N__19341\
        );

    \I__3160\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19341\
        );

    \I__3159\ : InMux
    port map (
            O => \N__19380\,
            I => \N__19341\
        );

    \I__3158\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19341\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19338\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19329\
        );

    \I__3155\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19329\
        );

    \I__3154\ : InMux
    port map (
            O => \N__19375\,
            I => \N__19329\
        );

    \I__3153\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19329\
        );

    \I__3152\ : InMux
    port map (
            O => \N__19373\,
            I => \N__19316\
        );

    \I__3151\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19316\
        );

    \I__3150\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19316\
        );

    \I__3149\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19316\
        );

    \I__3148\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19316\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19313\
        );

    \I__3146\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19310\
        );

    \I__3145\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19307\
        );

    \I__3144\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19302\
        );

    \I__3143\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19302\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__19359\,
            I => \N__19291\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__19352\,
            I => \N__19291\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19284\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19284\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__19329\,
            I => \N__19284\
        );

    \I__3137\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19279\
        );

    \I__3136\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19279\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__19316\,
            I => \N__19276\
        );

    \I__3134\ : Span4Mux_h
    port map (
            O => \N__19313\,
            I => \N__19267\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__19310\,
            I => \N__19267\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__19307\,
            I => \N__19267\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__19302\,
            I => \N__19267\
        );

    \I__3130\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19253\
        );

    \I__3129\ : InMux
    port map (
            O => \N__19300\,
            I => \N__19253\
        );

    \I__3128\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19253\
        );

    \I__3127\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19253\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19253\
        );

    \I__3125\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19253\
        );

    \I__3124\ : Span4Mux_s2_v
    port map (
            O => \N__19291\,
            I => \N__19250\
        );

    \I__3123\ : Span4Mux_v
    port map (
            O => \N__19284\,
            I => \N__19241\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__19279\,
            I => \N__19241\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__19276\,
            I => \N__19241\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__19267\,
            I => \N__19241\
        );

    \I__3119\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19238\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__19253\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__3117\ : Odrv4
    port map (
            O => \N__19250\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__19241\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19238\,
            I => \M_this_oam_ram_write_data_0_sqmuxa\
        );

    \I__3114\ : InMux
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19223\
        );

    \I__3112\ : Span4Mux_s3_v
    port map (
            O => \N__19223\,
            I => \N__19220\
        );

    \I__3111\ : Span4Mux_h
    port map (
            O => \N__19220\,
            I => \N__19217\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__19217\,
            I => \M_this_oam_ram_write_data_0\
        );

    \I__3109\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__19211\,
            I => \M_this_data_tmp_qZ0Z_0\
        );

    \I__3107\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19205\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__19205\,
            I => \M_this_data_tmp_qZ0Z_4\
        );

    \I__3105\ : InMux
    port map (
            O => \N__19202\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_6\
        );

    \I__3104\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__19196\,
            I => \this_ppu.M_state_q_RNISP3R6_1Z0Z_10\
        );

    \I__3102\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__3100\ : Span12Mux_h
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__3099\ : Odrv12
    port map (
            O => \N__19184\,
            I => \M_this_oam_ram_read_data_11\
        );

    \I__3098\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__3096\ : Span4Mux_v
    port map (
            O => \N__19175\,
            I => \N__19172\
        );

    \I__3095\ : Span4Mux_h
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__3094\ : Odrv4
    port map (
            O => \N__19169\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_11\
        );

    \I__3093\ : InMux
    port map (
            O => \N__19166\,
            I => \N__19163\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__19163\,
            I => \this_ppu.M_state_q_RNISP3R6Z0Z_10\
        );

    \I__3091\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19152\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19149\
        );

    \I__3089\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19140\
        );

    \I__3088\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19140\
        );

    \I__3087\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19140\
        );

    \I__3086\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19140\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__19152\,
            I => \this_ppu.N_806\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__19149\,
            I => \this_ppu.N_806\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__19140\,
            I => \this_ppu.N_806\
        );

    \I__3082\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19130\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__19130\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1\
        );

    \I__3080\ : InMux
    port map (
            O => \N__19127\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_0\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19124\,
            I => \N__19121\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__19121\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2\
        );

    \I__3077\ : InMux
    port map (
            O => \N__19118\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_1\
        );

    \I__3076\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19111\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19114\,
            I => \N__19108\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__19111\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_3\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__19108\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_3\
        );

    \I__3072\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19100\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__19100\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3\
        );

    \I__3070\ : InMux
    port map (
            O => \N__19097\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_2\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__19094\,
            I => \N__19091\
        );

    \I__3068\ : InMux
    port map (
            O => \N__19091\,
            I => \N__19087\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19090\,
            I => \N__19084\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__19087\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_4\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__19084\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_4\
        );

    \I__3064\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19076\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__19076\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4\
        );

    \I__3062\ : InMux
    port map (
            O => \N__19073\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_3\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19063\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19060\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19063\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_5\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__19060\,
            I => \this_ppu.M_pixel_cnt_qZ1Z_5\
        );

    \I__3056\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__19052\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5\
        );

    \I__3054\ : InMux
    port map (
            O => \N__19049\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_4\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__3052\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19039\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__19042\,
            I => \N__19036\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__19039\,
            I => \N__19033\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__19033\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_6\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19030\,
            I => \this_ppu.M_pixel_cnt_qZ0Z_6\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19022\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__3044\ : Span4Mux_h
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__19016\,
            I => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6\
        );

    \I__3042\ : InMux
    port map (
            O => \N__19013\,
            I => \this_ppu.un1_M_pixel_cnt_q_1_cry_5\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__19010\,
            I => \this_ppu.m9_0_a2_5_cascade_\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19007\,
            I => \N__19004\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__19004\,
            I => \this_vga_signals.i22_mux\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18997\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18993\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__18997\,
            I => \N__18990\
        );

    \I__3035\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18987\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__18993\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__3033\ : Odrv4
    port map (
            O => \N__18990\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__18987\,
            I => \this_vga_signals.M_lcounter_qZ0Z_1\
        );

    \I__3031\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18971\
        );

    \I__3030\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18971\
        );

    \I__3029\ : InMux
    port map (
            O => \N__18978\,
            I => \N__18971\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__18971\,
            I => \this_vga_signals.M_lcounter_qZ0Z_0\
        );

    \I__3027\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__18965\,
            I => \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__18962\,
            I => \this_ppu.N_814_cascade_\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__18959\,
            I => \this_ppu.N_806_cascade_\
        );

    \I__3023\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18950\
        );

    \I__3022\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18950\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__18950\,
            I => \this_ppu.un1_M_oam_curr_q_1_c5\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__3019\ : CascadeBuf
    port map (
            O => \N__18944\,
            I => \N__18941\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18938\
        );

    \I__3017\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__18935\,
            I => \N__18932\
        );

    \I__3015\ : Span4Mux_h
    port map (
            O => \N__18932\,
            I => \N__18929\
        );

    \I__3014\ : Span4Mux_v
    port map (
            O => \N__18929\,
            I => \N__18923\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__18928\,
            I => \N__18920\
        );

    \I__3012\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18917\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__18926\,
            I => \N__18914\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__18923\,
            I => \N__18911\
        );

    \I__3009\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18908\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__18917\,
            I => \N__18905\
        );

    \I__3007\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18902\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__18911\,
            I => \N__18899\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__18908\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__18905\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__18902\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__18899\,
            I => \M_this_ppu_oam_addr_5\
        );

    \I__3001\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18882\
        );

    \I__3000\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18877\
        );

    \I__2999\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18877\
        );

    \I__2998\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18874\
        );

    \I__2997\ : InMux
    port map (
            O => \N__18886\,
            I => \N__18869\
        );

    \I__2996\ : InMux
    port map (
            O => \N__18885\,
            I => \N__18869\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__18882\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__18877\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__18874\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__18869\,
            I => \this_ppu.M_oam_curr_qc_0_1\
        );

    \I__2991\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18856\
        );

    \I__2990\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18853\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__18853\,
            I => \this_ppu.M_oam_curr_qZ0Z_6\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__18850\,
            I => \this_ppu.M_oam_curr_qZ0Z_6\
        );

    \I__2986\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18838\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__18838\,
            I => \N__18832\
        );

    \I__2982\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18828\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__18832\,
            I => \N__18825\
        );

    \I__2980\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18822\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__18828\,
            I => \N__18819\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__18825\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__18822\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__2976\ : Odrv12
    port map (
            O => \N__18819\,
            I => \M_this_status_flags_qZ0Z_0\
        );

    \I__2975\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__18803\,
            I => \this_ppu.oam_cache.mem_15\
        );

    \I__2971\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18791\
        );

    \I__2970\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18791\
        );

    \I__2969\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18791\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__18788\,
            I => \N__18784\
        );

    \I__2966\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18781\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__18784\,
            I => \this_ppu.N_784_0\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__18781\,
            I => \this_ppu.N_784_0\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \this_vga_signals.N_859_cascade_\
        );

    \I__2962\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18770\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__18770\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_13\
        );

    \I__2960\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18764\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__18764\,
            I => \this_spr_ram.mem_mem_3_1_RNISI5GZ0\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__18761\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\
        );

    \I__2957\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18755\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__18755\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__18752\,
            I => \N__18749\
        );

    \I__2954\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18743\
        );

    \I__2953\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18740\
        );

    \I__2952\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18737\
        );

    \I__2951\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18734\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__18743\,
            I => \N__18731\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18726\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18726\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__18734\,
            I => \N__18723\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__18731\,
            I => \N__18718\
        );

    \I__2945\ : Span4Mux_v
    port map (
            O => \N__18726\,
            I => \N__18718\
        );

    \I__2944\ : Span4Mux_v
    port map (
            O => \N__18723\,
            I => \N__18713\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__18718\,
            I => \N__18713\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__18713\,
            I => \this_ppu_N_247\
        );

    \I__2941\ : InMux
    port map (
            O => \N__18710\,
            I => \N__18707\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__18707\,
            I => \N__18703\
        );

    \I__2939\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18700\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__18703\,
            I => \this_vga_signals.N_22_0\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__18700\,
            I => \this_vga_signals.N_22_0\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__18695\,
            I => \M_this_spr_ram_read_data_2_cascade_\
        );

    \I__2935\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18689\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__18689\,
            I => \N__18686\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__18686\,
            I => \N__18683\
        );

    \I__2932\ : Odrv4
    port map (
            O => \N__18683\,
            I => \N_28_0_i\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__18680\,
            I => \N__18677\
        );

    \I__2930\ : CascadeBuf
    port map (
            O => \N__18677\,
            I => \N__18674\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__18674\,
            I => \N__18671\
        );

    \I__2928\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18667\
        );

    \I__2927\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18663\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18660\
        );

    \I__2925\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18657\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__18663\,
            I => \N__18654\
        );

    \I__2923\ : Span4Mux_h
    port map (
            O => \N__18660\,
            I => \N__18651\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__18657\,
            I => \N__18647\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__18654\,
            I => \N__18643\
        );

    \I__2920\ : Sp12to4
    port map (
            O => \N__18651\,
            I => \N__18640\
        );

    \I__2919\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18637\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__18647\,
            I => \N__18634\
        );

    \I__2917\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18631\
        );

    \I__2916\ : Sp12to4
    port map (
            O => \N__18643\,
            I => \N__18626\
        );

    \I__2915\ : Span12Mux_s7_v
    port map (
            O => \N__18640\,
            I => \N__18626\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__18637\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__2913\ : Odrv4
    port map (
            O => \N__18634\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__18631\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__2911\ : Odrv12
    port map (
            O => \N__18626\,
            I => \M_this_ppu_oam_addr_4\
        );

    \I__2910\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__18614\,
            I => \M_this_spr_ram_read_data_2\
        );

    \I__2908\ : InMux
    port map (
            O => \N__18611\,
            I => \N__18607\
        );

    \I__2907\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18604\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__18607\,
            I => \N__18599\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__18604\,
            I => \N__18599\
        );

    \I__2904\ : Odrv12
    port map (
            O => \N__18599\,
            I => \M_this_spr_ram_read_data_1\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__2902\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__2899\ : Odrv4
    port map (
            O => \N__18584\,
            I => \M_this_spr_ram_read_data_3\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__18581\,
            I => \this_ppu.M_oam_curr_dZ0Z25_cascade_\
        );

    \I__2897\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__18572\,
            I => \N__18567\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18564\
        );

    \I__2893\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18561\
        );

    \I__2892\ : Span4Mux_v
    port map (
            O => \N__18567\,
            I => \N__18558\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__18564\,
            I => \this_ppu.N_834_0\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__18561\,
            I => \this_ppu.N_834_0\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__18558\,
            I => \this_ppu.N_834_0\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__2887\ : CascadeBuf
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__18545\,
            I => \N__18541\
        );

    \I__2885\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18537\
        );

    \I__2884\ : InMux
    port map (
            O => \N__18541\,
            I => \N__18534\
        );

    \I__2883\ : InMux
    port map (
            O => \N__18540\,
            I => \N__18530\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__18537\,
            I => \N__18527\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__18534\,
            I => \N__18524\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18521\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__18530\,
            I => \N__18518\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__18527\,
            I => \N__18514\
        );

    \I__2877\ : Span12Mux_s10_h
    port map (
            O => \N__18524\,
            I => \N__18510\
        );

    \I__2876\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18507\
        );

    \I__2875\ : Span4Mux_v
    port map (
            O => \N__18518\,
            I => \N__18504\
        );

    \I__2874\ : InMux
    port map (
            O => \N__18517\,
            I => \N__18501\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__18514\,
            I => \N__18498\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18495\
        );

    \I__2871\ : Span12Mux_v
    port map (
            O => \N__18510\,
            I => \N__18492\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__18507\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__18504\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__18501\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2867\ : Odrv4
    port map (
            O => \N__18498\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__18495\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2865\ : Odrv12
    port map (
            O => \N__18492\,
            I => \M_this_ppu_oam_addr_0\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__18479\,
            I => \this_ppu.N_834_0_cascade_\
        );

    \I__2863\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18472\
        );

    \I__2862\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18469\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__18472\,
            I => \N__18463\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__18469\,
            I => \N__18463\
        );

    \I__2859\ : InMux
    port map (
            O => \N__18468\,
            I => \N__18460\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__18460\,
            I => \this_ppu.un1_M_state_q_7_i_0_0\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__18457\,
            I => \this_ppu.un1_M_state_q_7_i_0_0\
        );

    \I__2855\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18446\
        );

    \I__2854\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18446\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18441\
        );

    \I__2852\ : InMux
    port map (
            O => \N__18445\,
            I => \N__18438\
        );

    \I__2851\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18435\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__18441\,
            I => \N__18432\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__18438\,
            I => \this_ppu.un1_M_oam_curr_q_1_c1\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__18435\,
            I => \this_ppu.un1_M_oam_curr_q_1_c1\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__18432\,
            I => \this_ppu.un1_M_oam_curr_q_1_c1\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__18425\,
            I => \N__18422\
        );

    \I__2845\ : CascadeBuf
    port map (
            O => \N__18422\,
            I => \N__18419\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__2843\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__2841\ : Span4Mux_v
    port map (
            O => \N__18410\,
            I => \N__18404\
        );

    \I__2840\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18399\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18399\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18396\
        );

    \I__2837\ : Sp12to4
    port map (
            O => \N__18404\,
            I => \N__18393\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__18399\,
            I => \N__18389\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__18396\,
            I => \N__18381\
        );

    \I__2834\ : Span12Mux_s6_h
    port map (
            O => \N__18393\,
            I => \N__18381\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18392\,
            I => \N__18378\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__18389\,
            I => \N__18375\
        );

    \I__2831\ : InMux
    port map (
            O => \N__18388\,
            I => \N__18370\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18370\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18367\
        );

    \I__2828\ : Span12Mux_v
    port map (
            O => \N__18381\,
            I => \N__18364\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__18378\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__18375\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__18370\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__18367\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__18364\,
            I => \M_this_ppu_oam_addr_1\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__18353\,
            I => \this_ppu.un1_M_oam_curr_q_1_c1_cascade_\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__18350\,
            I => \N__18346\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__18349\,
            I => \N__18343\
        );

    \I__2819\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18340\
        );

    \I__2818\ : CascadeBuf
    port map (
            O => \N__18343\,
            I => \N__18336\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__18340\,
            I => \N__18333\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18330\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__18336\,
            I => \N__18327\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__18333\,
            I => \N__18324\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18321\
        );

    \I__2812\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__2811\ : Sp12to4
    port map (
            O => \N__18324\,
            I => \N__18314\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__18321\,
            I => \N__18311\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__18318\,
            I => \N__18308\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__18317\,
            I => \N__18305\
        );

    \I__2807\ : Span12Mux_h
    port map (
            O => \N__18314\,
            I => \N__18296\
        );

    \I__2806\ : Sp12to4
    port map (
            O => \N__18311\,
            I => \N__18296\
        );

    \I__2805\ : Span12Mux_s10_h
    port map (
            O => \N__18308\,
            I => \N__18296\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18293\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18290\
        );

    \I__2802\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18287\
        );

    \I__2801\ : Span12Mux_v
    port map (
            O => \N__18296\,
            I => \N__18284\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__18293\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18290\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18287\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__2797\ : Odrv12
    port map (
            O => \N__18284\,
            I => \M_this_ppu_oam_addr_2\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18268\
        );

    \I__2795\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18265\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__18268\,
            I => \this_ppu.un1_M_oam_curr_q_1_c3\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__18265\,
            I => \this_ppu.un1_M_oam_curr_q_1_c3\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__2790\ : CascadeBuf
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__2788\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18248\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__18248\,
            I => \N__18244\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__18244\,
            I => \N__18237\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__18241\,
            I => \N__18233\
        );

    \I__2783\ : InMux
    port map (
            O => \N__18240\,
            I => \N__18230\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__18237\,
            I => \N__18227\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18224\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__18233\,
            I => \N__18218\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__18230\,
            I => \N__18213\
        );

    \I__2778\ : Span4Mux_v
    port map (
            O => \N__18227\,
            I => \N__18213\
        );

    \I__2777\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18208\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18208\
        );

    \I__2775\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18203\
        );

    \I__2774\ : InMux
    port map (
            O => \N__18221\,
            I => \N__18203\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__18218\,
            I => \N__18200\
        );

    \I__2772\ : Span4Mux_v
    port map (
            O => \N__18213\,
            I => \N__18197\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__18208\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__18203\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__18200\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__18197\,
            I => \M_this_ppu_oam_addr_3\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \this_ppu.un1_M_oam_curr_q_1_c3_cascade_\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__18185\,
            I => \N__18182\
        );

    \I__2765\ : CascadeBuf
    port map (
            O => \N__18182\,
            I => \N__18179\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__18179\,
            I => \N__18176\
        );

    \I__2763\ : InMux
    port map (
            O => \N__18176\,
            I => \N__18173\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__18173\,
            I => \N__18170\
        );

    \I__2761\ : Span4Mux_v
    port map (
            O => \N__18170\,
            I => \N__18167\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__18164\,
            I => \this_ppu.N_778_0\
        );

    \I__2758\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__18158\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_14\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__18152\,
            I => \N__18149\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__18149\,
            I => \N__18146\
        );

    \I__2753\ : Span4Mux_h
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__2752\ : Sp12to4
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__2751\ : Odrv12
    port map (
            O => \N__18140\,
            I => \this_spr_ram.mem_out_bus4_2\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18134\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__18134\,
            I => \N__18131\
        );

    \I__2748\ : Span12Mux_v
    port map (
            O => \N__18131\,
            I => \N__18128\
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__18128\,
            I => \this_spr_ram.mem_out_bus0_2\
        );

    \I__2746\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18122\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18122\,
            I => \N__18119\
        );

    \I__2744\ : Span4Mux_h
    port map (
            O => \N__18119\,
            I => \N__18116\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__18116\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_6\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__18113\,
            I => \this_ppu.M_state_q_inv_1_cascade_\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18107\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__18107\,
            I => \N__18104\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__18104\,
            I => \N__18101\
        );

    \I__2738\ : Sp12to4
    port map (
            O => \N__18101\,
            I => \N__18098\
        );

    \I__2737\ : Span12Mux_h
    port map (
            O => \N__18098\,
            I => \N__18095\
        );

    \I__2736\ : Span12Mux_v
    port map (
            O => \N__18095\,
            I => \N__18092\
        );

    \I__2735\ : Odrv12
    port map (
            O => \N__18092\,
            I => \M_this_map_ram_read_data_6\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__18089\,
            I => \N__18086\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18083\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__18083\,
            I => \N__18080\
        );

    \I__2731\ : Odrv12
    port map (
            O => \N__18080\,
            I => \this_ppu.m48_i_a2_0\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18074\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__18074\,
            I => \N__18071\
        );

    \I__2728\ : Span4Mux_v
    port map (
            O => \N__18071\,
            I => \N__18068\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__18068\,
            I => \N__18065\
        );

    \I__2726\ : Sp12to4
    port map (
            O => \N__18065\,
            I => \N__18062\
        );

    \I__2725\ : Odrv12
    port map (
            O => \N__18062\,
            I => \this_spr_ram.mem_out_bus5_2\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18056\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__2722\ : Span12Mux_v
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__2721\ : Span12Mux_v
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__2720\ : Odrv12
    port map (
            O => \N__18047\,
            I => \this_spr_ram.mem_out_bus1_2\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18044\,
            I => \N__18041\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__2717\ : Sp12to4
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__2716\ : Span12Mux_v
    port map (
            O => \N__18035\,
            I => \N__18032\
        );

    \I__2715\ : Odrv12
    port map (
            O => \N__18032\,
            I => \this_spr_ram.mem_out_bus7_2\
        );

    \I__2714\ : InMux
    port map (
            O => \N__18029\,
            I => \N__18026\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__18023\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__18023\,
            I => \N__18020\
        );

    \I__2711\ : Sp12to4
    port map (
            O => \N__18020\,
            I => \N__18017\
        );

    \I__2710\ : Span12Mux_h
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__18014\,
            I => \this_spr_ram.mem_out_bus3_2\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__2706\ : Sp12to4
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__2705\ : Span12Mux_v
    port map (
            O => \N__18002\,
            I => \N__17999\
        );

    \I__2704\ : Span12Mux_h
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__2703\ : Odrv12
    port map (
            O => \N__17996\,
            I => \this_spr_ram.mem_out_bus2_2\
        );

    \I__2702\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17990\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__2700\ : Span12Mux_v
    port map (
            O => \N__17987\,
            I => \N__17984\
        );

    \I__2699\ : Odrv12
    port map (
            O => \N__17984\,
            I => \this_spr_ram.mem_out_bus6_2\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__17981\,
            I => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_\
        );

    \I__2697\ : InMux
    port map (
            O => \N__17978\,
            I => \N__17975\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__17975\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\
        );

    \I__2695\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17969\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__17969\,
            I => \N__17966\
        );

    \I__2693\ : Sp12to4
    port map (
            O => \N__17966\,
            I => \N__17963\
        );

    \I__2692\ : Span12Mux_v
    port map (
            O => \N__17963\,
            I => \N__17960\
        );

    \I__2691\ : Span12Mux_h
    port map (
            O => \N__17960\,
            I => \N__17957\
        );

    \I__2690\ : Odrv12
    port map (
            O => \N__17957\,
            I => \this_spr_ram.mem_out_bus6_1\
        );

    \I__2689\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17951\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__17951\,
            I => \N__17948\
        );

    \I__2687\ : Sp12to4
    port map (
            O => \N__17948\,
            I => \N__17945\
        );

    \I__2686\ : Span12Mux_v
    port map (
            O => \N__17945\,
            I => \N__17942\
        );

    \I__2685\ : Span12Mux_h
    port map (
            O => \N__17942\,
            I => \N__17939\
        );

    \I__2684\ : Odrv12
    port map (
            O => \N__17939\,
            I => \this_spr_ram.mem_out_bus2_1\
        );

    \I__2683\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__17933\,
            I => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\
        );

    \I__2681\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17927\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__17927\,
            I => \N__17924\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__17924\,
            I => \N__17921\
        );

    \I__2678\ : Sp12to4
    port map (
            O => \N__17921\,
            I => \N__17918\
        );

    \I__2677\ : Odrv12
    port map (
            O => \N__17918\,
            I => \this_spr_ram.mem_out_bus4_3\
        );

    \I__2676\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17909\
        );

    \I__2674\ : Span12Mux_v
    port map (
            O => \N__17909\,
            I => \N__17906\
        );

    \I__2673\ : Odrv12
    port map (
            O => \N__17906\,
            I => \this_spr_ram.mem_out_bus0_3\
        );

    \I__2672\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17900\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__17900\,
            I => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__17897\,
            I => \N__17893\
        );

    \I__2669\ : InMux
    port map (
            O => \N__17896\,
            I => \N__17889\
        );

    \I__2668\ : InMux
    port map (
            O => \N__17893\,
            I => \N__17886\
        );

    \I__2667\ : InMux
    port map (
            O => \N__17892\,
            I => \N__17881\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17877\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__17886\,
            I => \N__17874\
        );

    \I__2664\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17869\
        );

    \I__2663\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17869\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__17881\,
            I => \N__17866\
        );

    \I__2661\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17863\
        );

    \I__2660\ : Span4Mux_v
    port map (
            O => \N__17877\,
            I => \N__17860\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__17874\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__17869\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__2657\ : Odrv12
    port map (
            O => \N__17866\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__17863\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__17860\,
            I => \M_this_ppu_vram_addr_3\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__17849\,
            I => \this_vga_signals.N_22_0_cascade_\
        );

    \I__2653\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__2651\ : Span4Mux_h
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__2650\ : Span4Mux_v
    port map (
            O => \N__17837\,
            I => \N__17834\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__17834\,
            I => \N_856_i\
        );

    \I__2648\ : InMux
    port map (
            O => \N__17831\,
            I => \N__17828\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__17828\,
            I => \N__17825\
        );

    \I__2646\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17822\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__2644\ : Sp12to4
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__2643\ : Odrv12
    port map (
            O => \N__17816\,
            I => \this_spr_ram.mem_out_bus5_3\
        );

    \I__2642\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17810\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__2640\ : Span12Mux_h
    port map (
            O => \N__17807\,
            I => \N__17804\
        );

    \I__2639\ : Span12Mux_v
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__2638\ : Odrv12
    port map (
            O => \N__17801\,
            I => \this_spr_ram.mem_out_bus1_3\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__17798\,
            I => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_\
        );

    \I__2636\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__17792\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__17789\,
            I => \M_this_spr_ram_read_data_3_cascade_\
        );

    \I__2633\ : InMux
    port map (
            O => \N__17786\,
            I => \N__17783\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__2631\ : Span12Mux_s11_h
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__2630\ : Odrv12
    port map (
            O => \N__17777\,
            I => \N_25_0_i\
        );

    \I__2629\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17771\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__17771\,
            I => \M_this_data_tmp_qZ0Z_23\
        );

    \I__2627\ : InMux
    port map (
            O => \N__17768\,
            I => \N__17765\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__17765\,
            I => \N__17762\
        );

    \I__2625\ : Span4Mux_h
    port map (
            O => \N__17762\,
            I => \N__17759\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__17759\,
            I => \M_this_oam_ram_write_data_19\
        );

    \I__2623\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17753\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17750\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__17750\,
            I => \M_this_oam_ram_write_data_28\
        );

    \I__2620\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17744\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17741\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__17741\,
            I => \M_this_oam_ram_write_data_25\
        );

    \I__2617\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17735\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__17735\,
            I => \N__17732\
        );

    \I__2615\ : Span4Mux_h
    port map (
            O => \N__17732\,
            I => \N__17729\
        );

    \I__2614\ : Sp12to4
    port map (
            O => \N__17729\,
            I => \N__17726\
        );

    \I__2613\ : Odrv12
    port map (
            O => \N__17726\,
            I => \this_spr_ram.mem_out_bus4_1\
        );

    \I__2612\ : InMux
    port map (
            O => \N__17723\,
            I => \N__17720\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17717\
        );

    \I__2610\ : Span4Mux_h
    port map (
            O => \N__17717\,
            I => \N__17714\
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__17714\,
            I => \this_spr_ram.mem_out_bus0_1\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__17708\,
            I => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__17705\,
            I => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\
        );

    \I__2605\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__2603\ : Span4Mux_v
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__2602\ : Span4Mux_h
    port map (
            O => \N__17693\,
            I => \N__17690\
        );

    \I__2601\ : Sp12to4
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__2600\ : Odrv12
    port map (
            O => \N__17687\,
            I => \this_spr_ram.mem_out_bus5_1\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17681\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__2597\ : Span12Mux_v
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__17675\,
            I => \this_spr_ram.mem_out_bus1_1\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17669\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__17669\,
            I => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\
        );

    \I__2593\ : InMux
    port map (
            O => \N__17666\,
            I => \N__17663\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17660\
        );

    \I__2591\ : Span12Mux_v
    port map (
            O => \N__17660\,
            I => \N__17657\
        );

    \I__2590\ : Span12Mux_v
    port map (
            O => \N__17657\,
            I => \N__17654\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__17654\,
            I => \this_spr_ram.mem_out_bus7_1\
        );

    \I__2588\ : InMux
    port map (
            O => \N__17651\,
            I => \N__17648\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__17648\,
            I => \N__17645\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__2585\ : Sp12to4
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__2584\ : Span12Mux_h
    port map (
            O => \N__17639\,
            I => \N__17636\
        );

    \I__2583\ : Odrv12
    port map (
            O => \N__17636\,
            I => \this_spr_ram.mem_out_bus3_1\
        );

    \I__2582\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17630\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__17630\,
            I => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\
        );

    \I__2580\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17624\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17621\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__17621\,
            I => \N__17618\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__17618\,
            I => \M_this_oam_ram_write_data_1\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17612\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17609\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__17609\,
            I => \M_this_data_tmp_qZ0Z_20\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17606\,
            I => \N__17603\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__2571\ : Span4Mux_h
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__17597\,
            I => \M_this_oam_ram_write_data_20\
        );

    \I__2569\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__17585\,
            I => \M_this_oam_ram_write_data_2\
        );

    \I__2565\ : InMux
    port map (
            O => \N__17582\,
            I => \N__17579\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__17579\,
            I => \M_this_data_tmp_qZ0Z_9\
        );

    \I__2563\ : InMux
    port map (
            O => \N__17576\,
            I => \N__17573\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__17570\,
            I => \M_this_oam_ram_write_data_9\
        );

    \I__2560\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17564\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__17558\,
            I => \M_this_oam_ram_write_data_4\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__17552\,
            I => \M_this_data_tmp_qZ0Z_11\
        );

    \I__2554\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2552\ : Odrv12
    port map (
            O => \N__17543\,
            I => \M_this_oam_ram_write_data_11\
        );

    \I__2551\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__17537\,
            I => \N__17534\
        );

    \I__2549\ : Span4Mux_s2_v
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__17531\,
            I => \M_this_data_tmp_qZ0Z_17\
        );

    \I__2547\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17525\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__17525\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_9\
        );

    \I__2545\ : InMux
    port map (
            O => \N__17522\,
            I => \N__17519\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17516\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__2542\ : Sp12to4
    port map (
            O => \N__17513\,
            I => \N__17509\
        );

    \I__2541\ : InMux
    port map (
            O => \N__17512\,
            I => \N__17506\
        );

    \I__2540\ : Odrv12
    port map (
            O => \N__17509\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__17506\,
            I => \this_ppu.M_oam_cache_read_data_16\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__17501\,
            I => \N__17498\
        );

    \I__2537\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17494\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__17497\,
            I => \N__17491\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__17494\,
            I => \N__17486\
        );

    \I__2534\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17483\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__17490\,
            I => \N__17480\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__17489\,
            I => \N__17476\
        );

    \I__2531\ : Span4Mux_s0_v
    port map (
            O => \N__17486\,
            I => \N__17470\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__17483\,
            I => \N__17470\
        );

    \I__2529\ : InMux
    port map (
            O => \N__17480\,
            I => \N__17467\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__17479\,
            I => \N__17464\
        );

    \I__2527\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17459\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__17475\,
            I => \N__17456\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__17470\,
            I => \N__17450\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__17467\,
            I => \N__17450\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17464\,
            I => \N__17447\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__17463\,
            I => \N__17444\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__17462\,
            I => \N__17440\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__17459\,
            I => \N__17436\
        );

    \I__2519\ : InMux
    port map (
            O => \N__17456\,
            I => \N__17433\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__17455\,
            I => \N__17430\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__17450\,
            I => \N__17423\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17423\
        );

    \I__2515\ : InMux
    port map (
            O => \N__17444\,
            I => \N__17420\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__17443\,
            I => \N__17417\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17414\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__17439\,
            I => \N__17411\
        );

    \I__2511\ : Span4Mux_s0_v
    port map (
            O => \N__17436\,
            I => \N__17406\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17406\
        );

    \I__2509\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17403\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__17429\,
            I => \N__17400\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__17428\,
            I => \N__17397\
        );

    \I__2506\ : Span4Mux_v
    port map (
            O => \N__17423\,
            I => \N__17392\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17392\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17389\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17414\,
            I => \N__17386\
        );

    \I__2502\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17383\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__17406\,
            I => \N__17378\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17378\
        );

    \I__2499\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17375\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17371\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__17392\,
            I => \N__17366\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__17389\,
            I => \N__17366\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__17386\,
            I => \N__17363\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__17383\,
            I => \N__17360\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__17378\,
            I => \N__17355\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__17375\,
            I => \N__17355\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__17374\,
            I => \N__17352\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__17371\,
            I => \N__17347\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__17366\,
            I => \N__17344\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__17363\,
            I => \N__17339\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__17360\,
            I => \N__17339\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__17355\,
            I => \N__17336\
        );

    \I__2485\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17333\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__17351\,
            I => \N__17330\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__17350\,
            I => \N__17327\
        );

    \I__2482\ : Span12Mux_h
    port map (
            O => \N__17347\,
            I => \N__17324\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__17344\,
            I => \N__17321\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__17339\,
            I => \N__17318\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__17336\,
            I => \N__17315\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__17333\,
            I => \N__17312\
        );

    \I__2477\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17309\
        );

    \I__2476\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17306\
        );

    \I__2475\ : Span12Mux_v
    port map (
            O => \N__17324\,
            I => \N__17301\
        );

    \I__2474\ : Sp12to4
    port map (
            O => \N__17321\,
            I => \N__17301\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__17318\,
            I => \N__17298\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__17315\,
            I => \N__17295\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__17312\,
            I => \N__17288\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__17309\,
            I => \N__17288\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__17306\,
            I => \N__17288\
        );

    \I__2468\ : Span12Mux_h
    port map (
            O => \N__17301\,
            I => \N__17285\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__17298\,
            I => \N__17282\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__17295\,
            I => \N__17277\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__17288\,
            I => \N__17277\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__17285\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__17282\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__17277\,
            I => \M_this_ppu_spr_addr_3\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \N__17267\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17260\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17255\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__17260\,
            I => \N__17252\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17259\,
            I => \N__17247\
        );

    \I__2455\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17247\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__17255\,
            I => \N__17244\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__17252\,
            I => \N__17241\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__17247\,
            I => \N__17238\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__17244\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__17241\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__2449\ : Odrv12
    port map (
            O => \N__17238\,
            I => \this_ppu.M_state_qZ0Z_2\
        );

    \I__2448\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \N__17228\
        );

    \I__2447\ : CascadeBuf
    port map (
            O => \N__17228\,
            I => \N__17225\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__2445\ : InMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__2443\ : Span4Mux_h
    port map (
            O => \N__17216\,
            I => \N__17211\
        );

    \I__2442\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17206\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17206\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__17211\,
            I => \N__17203\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__17206\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__17203\,
            I => \M_this_oam_address_qZ0Z_6\
        );

    \I__2437\ : CascadeMux
    port map (
            O => \N__17198\,
            I => \N__17195\
        );

    \I__2436\ : CascadeBuf
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2434\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__2432\ : Span4Mux_s2_v
    port map (
            O => \N__17183\,
            I => \N__17179\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__17176\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__17173\,
            I => \M_this_oam_address_qZ0Z_7\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__17165\,
            I => \M_this_data_tmp_qZ0Z_12\
        );

    \I__2425\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__17159\,
            I => \N__17156\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__17156\,
            I => \M_this_data_tmp_qZ0Z_15\
        );

    \I__2422\ : InMux
    port map (
            O => \N__17153\,
            I => \N__17150\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__17150\,
            I => \N__17147\
        );

    \I__2420\ : Odrv4
    port map (
            O => \N__17147\,
            I => \M_this_data_tmp_qZ0Z_13\
        );

    \I__2419\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17138\
        );

    \I__2418\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17131\
        );

    \I__2417\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17131\
        );

    \I__2416\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17131\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__17138\,
            I => \this_ppu.N_1210_0\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__17131\,
            I => \this_ppu.N_1210_0\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__17123\,
            I => \this_ppu.un1_M_screen_x_q_c3\
        );

    \I__2411\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17117\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__2409\ : Odrv12
    port map (
            O => \N__17114\,
            I => \this_ppu.oam_cache.mem_13\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__17105\,
            I => \this_ppu.oam_cache.mem_12\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__17096\,
            I => \this_ppu.m13_0_a2_0_0\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__17093\,
            I => \this_ppu.N_844_cascade_\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17084\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17089\,
            I => \N__17084\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17084\,
            I => \N__17080\
        );

    \I__2398\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__17080\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__17077\,
            I => \this_ppu.M_state_qZ0Z_1\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17068\
        );

    \I__2394\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17065\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__17068\,
            I => \M_this_warmup_qZ0Z_1\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__17065\,
            I => \M_this_warmup_qZ0Z_1\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__17060\,
            I => \N__17055\
        );

    \I__2390\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17050\
        );

    \I__2389\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17050\
        );

    \I__2388\ : InMux
    port map (
            O => \N__17055\,
            I => \N__17047\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__17050\,
            I => \M_this_warmup_qZ0Z_0\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17047\,
            I => \M_this_warmup_qZ0Z_0\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__17042\,
            I => \this_ppu.N_827_0_cascade_\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__17039\,
            I => \this_ppu.un1_M_screen_x_q_c2_cascade_\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17033\,
            I => \this_ppu.un1_M_screen_x_q_c5\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__17030\,
            I => \this_ppu.un1_M_screen_x_q_c5_cascade_\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__17018\,
            I => \N__17013\
        );

    \I__2376\ : InMux
    port map (
            O => \N__17017\,
            I => \N__17008\
        );

    \I__2375\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17008\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__17013\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17008\,
            I => \M_this_ppu_vram_addr_5\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__2371\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__16994\,
            I => \N__16990\
        );

    \I__2368\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16987\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__16990\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__16987\,
            I => \M_this_ppu_vram_addr_6\
        );

    \I__2365\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__16979\,
            I => \this_ppu.un1_M_screen_x_q_c2\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__2362\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16970\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__16967\,
            I => \N__16961\
        );

    \I__2359\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16958\
        );

    \I__2358\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16953\
        );

    \I__2357\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16953\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__16961\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__16958\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__16953\,
            I => \M_this_ppu_vram_addr_1\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__16946\,
            I => \N__16943\
        );

    \I__2352\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16938\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__16942\,
            I => \N__16935\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__16941\,
            I => \N__16932\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__16938\,
            I => \N__16929\
        );

    \I__2348\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16922\
        );

    \I__2347\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16922\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__16929\,
            I => \N__16919\
        );

    \I__2345\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16916\
        );

    \I__2344\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16913\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__16922\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__16919\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__16916\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__16913\,
            I => \M_this_ppu_vram_addr_0\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__16904\,
            I => \N__16901\
        );

    \I__2338\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16897\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__16900\,
            I => \N__16893\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16890\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__16896\,
            I => \N__16887\
        );

    \I__2334\ : InMux
    port map (
            O => \N__16893\,
            I => \N__16884\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__16890\,
            I => \N__16880\
        );

    \I__2332\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16877\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__16884\,
            I => \N__16874\
        );

    \I__2330\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16871\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__16880\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__16877\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__16874\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__16871\,
            I => \M_this_ppu_vram_addr_2\
        );

    \I__2325\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16855\
        );

    \I__2324\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16855\
        );

    \I__2323\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16852\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__16855\,
            I => \this_ppu.N_827_0\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__16852\,
            I => \this_ppu.N_827_0\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__16847\,
            I => \this_ppu.un1_M_screen_x_q_c3_cascade_\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__2318\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16838\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__16835\,
            I => \N__16830\
        );

    \I__2315\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16827\
        );

    \I__2314\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16824\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__16830\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__16827\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__16824\,
            I => \M_this_ppu_vram_addr_4\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__16817\,
            I => \this_ppu.M_oam_curr_qc_0_1_cascade_\
        );

    \I__2309\ : InMux
    port map (
            O => \N__16814\,
            I => \N__16811\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__16811\,
            I => \N__16808\
        );

    \I__2307\ : Span4Mux_h
    port map (
            O => \N__16808\,
            I => \N__16805\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__16805\,
            I => \this_ppu.m35_i_a2_4\
        );

    \I__2305\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16799\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__16799\,
            I => \N__16796\
        );

    \I__2303\ : Span4Mux_s1_v
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__16793\,
            I => \M_this_oam_ram_write_data_21\
        );

    \I__2301\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__16787\,
            I => \N__16784\
        );

    \I__2299\ : Span4Mux_s1_v
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__16781\,
            I => \M_this_oam_ram_write_data_23\
        );

    \I__2297\ : CEMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16771\
        );

    \I__2295\ : CEMux
    port map (
            O => \N__16774\,
            I => \N__16768\
        );

    \I__2294\ : Span4Mux_s3_v
    port map (
            O => \N__16771\,
            I => \N__16763\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__16768\,
            I => \N__16763\
        );

    \I__2292\ : Span4Mux_h
    port map (
            O => \N__16763\,
            I => \N__16760\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__16760\,
            I => \this_spr_ram.mem_WE_12\
        );

    \I__2290\ : CEMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__16754\,
            I => \N__16750\
        );

    \I__2288\ : CEMux
    port map (
            O => \N__16753\,
            I => \N__16747\
        );

    \I__2287\ : Span4Mux_v
    port map (
            O => \N__16750\,
            I => \N__16742\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__16747\,
            I => \N__16742\
        );

    \I__2285\ : Span4Mux_h
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__16739\,
            I => \this_spr_ram.mem_WE_14\
        );

    \I__2283\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16733\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__16730\,
            I => \N__16727\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__2279\ : Odrv4
    port map (
            O => \N__16724\,
            I => \this_ppu.oam_cache.mem_5\
        );

    \I__2278\ : CEMux
    port map (
            O => \N__16721\,
            I => \N__16718\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__16718\,
            I => \N__16715\
        );

    \I__2276\ : Span4Mux_v
    port map (
            O => \N__16715\,
            I => \N__16711\
        );

    \I__2275\ : CEMux
    port map (
            O => \N__16714\,
            I => \N__16708\
        );

    \I__2274\ : Sp12to4
    port map (
            O => \N__16711\,
            I => \N__16703\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__16708\,
            I => \N__16703\
        );

    \I__2272\ : Span12Mux_h
    port map (
            O => \N__16703\,
            I => \N__16700\
        );

    \I__2271\ : Span12Mux_v
    port map (
            O => \N__16700\,
            I => \N__16697\
        );

    \I__2270\ : Odrv12
    port map (
            O => \N__16697\,
            I => \this_spr_ram.mem_WE_0\
        );

    \I__2269\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16691\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__16691\,
            I => \N__16688\
        );

    \I__2267\ : Span4Mux_v
    port map (
            O => \N__16688\,
            I => \N__16685\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__16685\,
            I => \N_34_i\
        );

    \I__2265\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16676\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__16670\,
            I => \this_ppu.oam_cache.mem_14\
        );

    \I__2260\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__16664\,
            I => \M_this_data_tmp_qZ0Z_8\
        );

    \I__2258\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__16658\,
            I => \M_this_data_tmp_qZ0Z_14\
        );

    \I__2256\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16652\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__16652\,
            I => \M_this_data_tmp_qZ0Z_10\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__16643\,
            I => \N__16640\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__16640\,
            I => \M_this_oam_ram_write_data_10\
        );

    \I__2250\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__16628\,
            I => \M_this_oam_ram_write_data_12\
        );

    \I__2246\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__16622\,
            I => \M_this_data_tmp_qZ0Z_7\
        );

    \I__2244\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__16616\,
            I => \M_this_data_tmp_qZ0Z_5\
        );

    \I__2242\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__16610\,
            I => \M_this_data_tmp_qZ0Z_22\
        );

    \I__2240\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16604\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__16604\,
            I => \M_this_data_tmp_qZ0Z_16\
        );

    \I__2238\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__2236\ : Odrv4
    port map (
            O => \N__16595\,
            I => \M_this_oam_ram_write_data_31\
        );

    \I__2235\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__16589\,
            I => \M_this_warmup_qZ0Z_22\
        );

    \I__2233\ : InMux
    port map (
            O => \N__16586\,
            I => \un1_M_this_warmup_d_cry_21\
        );

    \I__2232\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16580\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__16580\,
            I => \M_this_warmup_qZ0Z_23\
        );

    \I__2230\ : InMux
    port map (
            O => \N__16577\,
            I => \un1_M_this_warmup_d_cry_22\
        );

    \I__2229\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__16571\,
            I => \M_this_warmup_qZ0Z_24\
        );

    \I__2227\ : InMux
    port map (
            O => \N__16568\,
            I => \un1_M_this_warmup_d_cry_23\
        );

    \I__2226\ : InMux
    port map (
            O => \N__16565\,
            I => \N__16562\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__16562\,
            I => \M_this_warmup_qZ0Z_25\
        );

    \I__2224\ : InMux
    port map (
            O => \N__16559\,
            I => \bfn_10_23_0_\
        );

    \I__2223\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__16553\,
            I => \M_this_warmup_qZ0Z_26\
        );

    \I__2221\ : InMux
    port map (
            O => \N__16550\,
            I => \un1_M_this_warmup_d_cry_25\
        );

    \I__2220\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__16544\,
            I => \M_this_warmup_qZ0Z_27\
        );

    \I__2218\ : InMux
    port map (
            O => \N__16541\,
            I => \un1_M_this_warmup_d_cry_26\
        );

    \I__2217\ : InMux
    port map (
            O => \N__16538\,
            I => \un1_M_this_warmup_d_cry_27\
        );

    \I__2216\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16529\
        );

    \I__2215\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16529\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__16529\,
            I => \M_this_warmup_qZ0Z_28\
        );

    \I__2213\ : InMux
    port map (
            O => \N__16526\,
            I => \un1_M_this_warmup_d_cry_12\
        );

    \I__2212\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__16520\,
            I => \M_this_warmup_qZ0Z_14\
        );

    \I__2210\ : InMux
    port map (
            O => \N__16517\,
            I => \un1_M_this_warmup_d_cry_13\
        );

    \I__2209\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__16511\,
            I => \M_this_warmup_qZ0Z_15\
        );

    \I__2207\ : InMux
    port map (
            O => \N__16508\,
            I => \un1_M_this_warmup_d_cry_14\
        );

    \I__2206\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__16502\,
            I => \M_this_warmup_qZ0Z_16\
        );

    \I__2204\ : InMux
    port map (
            O => \N__16499\,
            I => \un1_M_this_warmup_d_cry_15\
        );

    \I__2203\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__16493\,
            I => \M_this_warmup_qZ0Z_17\
        );

    \I__2201\ : InMux
    port map (
            O => \N__16490\,
            I => \bfn_10_22_0_\
        );

    \I__2200\ : InMux
    port map (
            O => \N__16487\,
            I => \N__16484\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__16484\,
            I => \M_this_warmup_qZ0Z_18\
        );

    \I__2198\ : InMux
    port map (
            O => \N__16481\,
            I => \un1_M_this_warmup_d_cry_17\
        );

    \I__2197\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16475\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__16475\,
            I => \M_this_warmup_qZ0Z_19\
        );

    \I__2195\ : InMux
    port map (
            O => \N__16472\,
            I => \un1_M_this_warmup_d_cry_18\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16469\,
            I => \N__16466\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__16466\,
            I => \M_this_warmup_qZ0Z_20\
        );

    \I__2192\ : InMux
    port map (
            O => \N__16463\,
            I => \un1_M_this_warmup_d_cry_19\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__16457\,
            I => \M_this_warmup_qZ0Z_21\
        );

    \I__2189\ : InMux
    port map (
            O => \N__16454\,
            I => \un1_M_this_warmup_d_cry_20\
        );

    \I__2188\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__16448\,
            I => \M_this_warmup_qZ0Z_5\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16445\,
            I => \un1_M_this_warmup_d_cry_4\
        );

    \I__2185\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16439\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__16439\,
            I => \M_this_warmup_qZ0Z_6\
        );

    \I__2183\ : InMux
    port map (
            O => \N__16436\,
            I => \un1_M_this_warmup_d_cry_5\
        );

    \I__2182\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__16430\,
            I => \M_this_warmup_qZ0Z_7\
        );

    \I__2180\ : InMux
    port map (
            O => \N__16427\,
            I => \un1_M_this_warmup_d_cry_6\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__16421\,
            I => \M_this_warmup_qZ0Z_8\
        );

    \I__2177\ : InMux
    port map (
            O => \N__16418\,
            I => \un1_M_this_warmup_d_cry_7\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__16412\,
            I => \M_this_warmup_qZ0Z_9\
        );

    \I__2174\ : InMux
    port map (
            O => \N__16409\,
            I => \bfn_10_21_0_\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__16403\,
            I => \M_this_warmup_qZ0Z_10\
        );

    \I__2171\ : InMux
    port map (
            O => \N__16400\,
            I => \un1_M_this_warmup_d_cry_9\
        );

    \I__2170\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__16394\,
            I => \M_this_warmup_qZ0Z_11\
        );

    \I__2168\ : InMux
    port map (
            O => \N__16391\,
            I => \un1_M_this_warmup_d_cry_10\
        );

    \I__2167\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__16385\,
            I => \M_this_warmup_qZ0Z_12\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16382\,
            I => \un1_M_this_warmup_d_cry_11\
        );

    \I__2164\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16376\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__16376\,
            I => \M_this_warmup_qZ0Z_13\
        );

    \I__2162\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__16367\,
            I => \this_ppu.oam_cache.mem_10\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__16358\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_10\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__16355\,
            I => \this_ppu.N_836_cascade_\
        );

    \I__2155\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16349\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__16349\,
            I => \N__16346\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__16346\,
            I => \N__16343\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__16343\,
            I => \this_ppu.oam_cache.mem_9\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__16337\,
            I => \M_this_warmup_qZ0Z_2\
        );

    \I__2149\ : InMux
    port map (
            O => \N__16334\,
            I => \un1_M_this_warmup_d_cry_1\
        );

    \I__2148\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__16328\,
            I => \M_this_warmup_qZ0Z_3\
        );

    \I__2146\ : InMux
    port map (
            O => \N__16325\,
            I => \un1_M_this_warmup_d_cry_2\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16319\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__16319\,
            I => \M_this_warmup_qZ0Z_4\
        );

    \I__2143\ : InMux
    port map (
            O => \N__16316\,
            I => \un1_M_this_warmup_d_cry_3\
        );

    \I__2142\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16310\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__16310\,
            I => \N__16307\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__16307\,
            I => \N__16303\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__16303\,
            I => \this_vga_signals.M_pcounter_q_i_2_0\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__16300\,
            I => \this_vga_signals.M_pcounter_q_i_2_0\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16292\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__16292\,
            I => \this_vga_signals.M_pcounter_q_3_0\
        );

    \I__2134\ : SRMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__16286\,
            I => \N__16282\
        );

    \I__2132\ : SRMux
    port map (
            O => \N__16285\,
            I => \N__16279\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__16282\,
            I => \N__16275\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__16279\,
            I => \N__16272\
        );

    \I__2129\ : SRMux
    port map (
            O => \N__16278\,
            I => \N__16269\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__16275\,
            I => \this_vga_signals.N_1188_1\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__16272\,
            I => \this_vga_signals.N_1188_1\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__16269\,
            I => \this_vga_signals.N_1188_1\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__16262\,
            I => \this_vga_signals.N_1188_1_cascade_\
        );

    \I__2124\ : CEMux
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__16256\,
            I => \N__16253\
        );

    \I__2122\ : Span4Mux_h
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__16250\,
            I => \this_vga_signals.N_933_1\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16244\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16238\
        );

    \I__2118\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16235\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16232\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16229\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__16238\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__16235\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__16232\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__16229\,
            I => \this_vga_signals.M_pcounter_qZ0Z_1\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__16220\,
            I => \N__16216\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__16219\,
            I => \N__16212\
        );

    \I__2109\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16207\
        );

    \I__2108\ : InMux
    port map (
            O => \N__16215\,
            I => \N__16207\
        );

    \I__2107\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16204\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__16204\,
            I => \N__16196\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__16201\,
            I => \N__16196\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__16196\,
            I => \this_vga_signals.M_pcounter_qZ0Z_0\
        );

    \I__2102\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__16190\,
            I => \N_2_0\
        );

    \I__2100\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__16184\,
            I => \M_this_vga_signals_pixel_clk_0_0\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__16181\,
            I => \N_2_0_cascade_\
        );

    \I__2097\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16172\
        );

    \I__2096\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16172\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N_3_0\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__16166\,
            I => \N__16161\
        );

    \I__2092\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16152\
        );

    \I__2091\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16152\
        );

    \I__2090\ : Span4Mux_h
    port map (
            O => \N__16161\,
            I => \N__16149\
        );

    \I__2089\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16146\
        );

    \I__2088\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16139\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16139\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16139\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16136\
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__16149\,
            I => \G_462\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__16146\,
            I => \G_462\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__16139\,
            I => \G_462\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__16136\,
            I => \G_462\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__16127\,
            I => \N__16124\
        );

    \I__2079\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16121\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__16121\,
            I => \this_ppu.M_oam_cache_read_data_i_16\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__2076\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16112\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16112\,
            I => \this_ppu.M_oam_cache_read_data_i_17\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__16109\,
            I => \N__16105\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__16108\,
            I => \N__16102\
        );

    \I__2072\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16098\
        );

    \I__2071\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16095\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__16101\,
            I => \N__16092\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16083\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__16095\,
            I => \N__16083\
        );

    \I__2067\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16080\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16077\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \N__16074\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__16089\,
            I => \N__16069\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__16088\,
            I => \N__16066\
        );

    \I__2062\ : Span4Mux_s2_v
    port map (
            O => \N__16083\,
            I => \N__16060\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16060\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16077\,
            I => \N__16057\
        );

    \I__2059\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16054\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__16073\,
            I => \N__16051\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__16072\,
            I => \N__16048\
        );

    \I__2056\ : InMux
    port map (
            O => \N__16069\,
            I => \N__16043\
        );

    \I__2055\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16040\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__16065\,
            I => \N__16037\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__16060\,
            I => \N__16032\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16032\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__16054\,
            I => \N__16029\
        );

    \I__2050\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16026\
        );

    \I__2049\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16023\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__16047\,
            I => \N__16020\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__16046\,
            I => \N__16017\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16012\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__16040\,
            I => \N__16012\
        );

    \I__2044\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16009\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__16032\,
            I => \N__15999\
        );

    \I__2042\ : Span4Mux_h
    port map (
            O => \N__16029\,
            I => \N__15999\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__15999\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__16023\,
            I => \N__15996\
        );

    \I__2039\ : InMux
    port map (
            O => \N__16020\,
            I => \N__15993\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16017\,
            I => \N__15990\
        );

    \I__2037\ : Span4Mux_s2_v
    port map (
            O => \N__16012\,
            I => \N__15985\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__16009\,
            I => \N__15985\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__16008\,
            I => \N__15982\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__16007\,
            I => \N__15979\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__16006\,
            I => \N__15976\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__15999\,
            I => \N__15968\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__15996\,
            I => \N__15968\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15968\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15965\
        );

    \I__2028\ : Span4Mux_v
    port map (
            O => \N__15985\,
            I => \N__15962\
        );

    \I__2027\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15959\
        );

    \I__2026\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15956\
        );

    \I__2025\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15953\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__15975\,
            I => \N__15950\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__15968\,
            I => \N__15947\
        );

    \I__2022\ : Span12Mux_h
    port map (
            O => \N__15965\,
            I => \N__15940\
        );

    \I__2021\ : Sp12to4
    port map (
            O => \N__15962\,
            I => \N__15940\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__15959\,
            I => \N__15940\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__15956\,
            I => \N__15937\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15934\
        );

    \I__2017\ : InMux
    port map (
            O => \N__15950\,
            I => \N__15931\
        );

    \I__2016\ : Sp12to4
    port map (
            O => \N__15947\,
            I => \N__15928\
        );

    \I__2015\ : Span12Mux_h
    port map (
            O => \N__15940\,
            I => \N__15925\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__15937\,
            I => \N__15918\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__15934\,
            I => \N__15918\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__15931\,
            I => \N__15918\
        );

    \I__2011\ : Span12Mux_h
    port map (
            O => \N__15928\,
            I => \N__15913\
        );

    \I__2010\ : Span12Mux_v
    port map (
            O => \N__15925\,
            I => \N__15913\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__15918\,
            I => \N__15910\
        );

    \I__2008\ : Odrv12
    port map (
            O => \N__15913\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__15910\,
            I => \M_this_ppu_spr_addr_4\
        );

    \I__2006\ : InMux
    port map (
            O => \N__15905\,
            I => \this_ppu.offset_y_cry_0\
        );

    \I__2005\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__15899\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_18\
        );

    \I__2003\ : InMux
    port map (
            O => \N__15896\,
            I => \this_ppu.offset_y_cry_1\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__2001\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15884\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__15889\,
            I => \N__15881\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__15888\,
            I => \N__15877\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__15887\,
            I => \N__15874\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__15884\,
            I => \N__15869\
        );

    \I__1996\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15866\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \N__15863\
        );

    \I__1994\ : InMux
    port map (
            O => \N__15877\,
            I => \N__15860\
        );

    \I__1993\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15857\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__15873\,
            I => \N__15850\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__15872\,
            I => \N__15847\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__15869\,
            I => \N__15841\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15841\
        );

    \I__1988\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15838\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__15860\,
            I => \N__15834\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__15857\,
            I => \N__15831\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15828\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15823\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__15854\,
            I => \N__15819\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__15853\,
            I => \N__15816\
        );

    \I__1981\ : InMux
    port map (
            O => \N__15850\,
            I => \N__15813\
        );

    \I__1980\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15810\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__15846\,
            I => \N__15807\
        );

    \I__1978\ : Span4Mux_v
    port map (
            O => \N__15841\,
            I => \N__15802\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__15838\,
            I => \N__15802\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__15837\,
            I => \N__15799\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__15834\,
            I => \N__15796\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__15831\,
            I => \N__15793\
        );

    \I__1973\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15790\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__15827\,
            I => \N__15787\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__15826\,
            I => \N__15784\
        );

    \I__1970\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15781\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__15822\,
            I => \N__15778\
        );

    \I__1968\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15775\
        );

    \I__1967\ : InMux
    port map (
            O => \N__15816\,
            I => \N__15772\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__15813\,
            I => \N__15769\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__15810\,
            I => \N__15766\
        );

    \I__1964\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15763\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__15802\,
            I => \N__15760\
        );

    \I__1962\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15757\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__15796\,
            I => \N__15754\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__15793\,
            I => \N__15751\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__15790\,
            I => \N__15748\
        );

    \I__1958\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15745\
        );

    \I__1957\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15742\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__15781\,
            I => \N__15739\
        );

    \I__1955\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15736\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__15775\,
            I => \N__15733\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__15772\,
            I => \N__15730\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__15769\,
            I => \N__15727\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__15766\,
            I => \N__15724\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__15763\,
            I => \N__15721\
        );

    \I__1949\ : Sp12to4
    port map (
            O => \N__15760\,
            I => \N__15718\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__15757\,
            I => \N__15715\
        );

    \I__1947\ : Sp12to4
    port map (
            O => \N__15754\,
            I => \N__15708\
        );

    \I__1946\ : Sp12to4
    port map (
            O => \N__15751\,
            I => \N__15708\
        );

    \I__1945\ : Span12Mux_s10_h
    port map (
            O => \N__15748\,
            I => \N__15708\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15705\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__15742\,
            I => \N__15702\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__15739\,
            I => \N__15699\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__15736\,
            I => \N__15696\
        );

    \I__1940\ : Span12Mux_h
    port map (
            O => \N__15733\,
            I => \N__15693\
        );

    \I__1939\ : Span12Mux_s10_h
    port map (
            O => \N__15730\,
            I => \N__15690\
        );

    \I__1938\ : Sp12to4
    port map (
            O => \N__15727\,
            I => \N__15687\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__15724\,
            I => \N__15682\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__15721\,
            I => \N__15682\
        );

    \I__1935\ : Span12Mux_v
    port map (
            O => \N__15718\,
            I => \N__15677\
        );

    \I__1934\ : Span12Mux_s10_h
    port map (
            O => \N__15715\,
            I => \N__15677\
        );

    \I__1933\ : Span12Mux_h
    port map (
            O => \N__15708\,
            I => \N__15672\
        );

    \I__1932\ : Span12Mux_s9_h
    port map (
            O => \N__15705\,
            I => \N__15672\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__15702\,
            I => \N__15669\
        );

    \I__1930\ : Span4Mux_v
    port map (
            O => \N__15699\,
            I => \N__15664\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__15696\,
            I => \N__15664\
        );

    \I__1928\ : Span12Mux_v
    port map (
            O => \N__15693\,
            I => \N__15661\
        );

    \I__1927\ : Span12Mux_h
    port map (
            O => \N__15690\,
            I => \N__15654\
        );

    \I__1926\ : Span12Mux_s8_v
    port map (
            O => \N__15687\,
            I => \N__15654\
        );

    \I__1925\ : Sp12to4
    port map (
            O => \N__15682\,
            I => \N__15654\
        );

    \I__1924\ : Span12Mux_h
    port map (
            O => \N__15677\,
            I => \N__15647\
        );

    \I__1923\ : Span12Mux_v
    port map (
            O => \N__15672\,
            I => \N__15647\
        );

    \I__1922\ : Sp12to4
    port map (
            O => \N__15669\,
            I => \N__15647\
        );

    \I__1921\ : Span4Mux_v
    port map (
            O => \N__15664\,
            I => \N__15644\
        );

    \I__1920\ : Odrv12
    port map (
            O => \N__15661\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1919\ : Odrv12
    port map (
            O => \N__15654\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1918\ : Odrv12
    port map (
            O => \N__15647\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__15644\,
            I => \M_this_ppu_spr_addr_5\
        );

    \I__1916\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__1914\ : Span4Mux_h
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__1913\ : Sp12to4
    port map (
            O => \N__15626\,
            I => \N__15623\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__15623\,
            I => \this_ppu.oam_cache.mem_4\
        );

    \I__1911\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15614\
        );

    \I__1910\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15614\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__15614\,
            I => \this_pixel_clk_M_counter_q_i_1\
        );

    \I__1908\ : InMux
    port map (
            O => \N__15611\,
            I => \N__15606\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15601\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15601\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__15606\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__15601\,
            I => \this_pixel_clk_M_counter_q_0\
        );

    \I__1903\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15593\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__15593\,
            I => \N__15588\
        );

    \I__1901\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15585\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__15591\,
            I => \N__15578\
        );

    \I__1899\ : Sp12to4
    port map (
            O => \N__15588\,
            I => \N__15572\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__15585\,
            I => \N__15572\
        );

    \I__1897\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15569\
        );

    \I__1896\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15560\
        );

    \I__1895\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15560\
        );

    \I__1894\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15560\
        );

    \I__1893\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15560\
        );

    \I__1892\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15556\
        );

    \I__1891\ : Span12Mux_v
    port map (
            O => \N__15572\,
            I => \N__15549\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15549\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__15560\,
            I => \N__15549\
        );

    \I__1888\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15546\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__15556\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__15549\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__15546\,
            I => \this_vga_signals.M_hcounter_qZ0Z_1\
        );

    \I__1884\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15535\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__15535\,
            I => \N__15526\
        );

    \I__1881\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15523\
        );

    \I__1880\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15520\
        );

    \I__1879\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15514\
        );

    \I__1878\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15514\
        );

    \I__1877\ : Span12Mux_v
    port map (
            O => \N__15526\,
            I => \N__15507\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__15523\,
            I => \N__15507\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__15520\,
            I => \N__15507\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15504\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15514\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__15507\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__15504\,
            I => \this_vga_signals.M_hcounter_qZ0Z_0\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__15497\,
            I => \N_3_0_cascade_\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15488\
        );

    \I__1868\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15488\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__15485\,
            I => \M_this_oam_ram_read_data_20\
        );

    \I__1865\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__1863\ : Span12Mux_v
    port map (
            O => \N__15476\,
            I => \N__15473\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__15473\,
            I => \M_this_oam_ram_read_data_i_20\
        );

    \I__1861\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__15467\,
            I => \M_this_oam_ram_write_data_27\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15461\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__15461\,
            I => \M_this_oam_ram_write_data_30\
        );

    \I__1857\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15455\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__15455\,
            I => \M_this_oam_ram_write_data_17\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__15449\,
            I => \M_this_oam_ram_write_data_29\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__15443\,
            I => \M_this_oam_ram_write_data_24\
        );

    \I__1851\ : IoInMux
    port map (
            O => \N__15440\,
            I => \N__15437\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__15437\,
            I => \N__15432\
        );

    \I__1849\ : IoInMux
    port map (
            O => \N__15436\,
            I => \N__15429\
        );

    \I__1848\ : IoInMux
    port map (
            O => \N__15435\,
            I => \N__15426\
        );

    \I__1847\ : IoSpan4Mux
    port map (
            O => \N__15432\,
            I => \N__15416\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__15429\,
            I => \N__15416\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__15426\,
            I => \N__15416\
        );

    \I__1844\ : IoInMux
    port map (
            O => \N__15425\,
            I => \N__15413\
        );

    \I__1843\ : IoInMux
    port map (
            O => \N__15424\,
            I => \N__15410\
        );

    \I__1842\ : IoInMux
    port map (
            O => \N__15423\,
            I => \N__15405\
        );

    \I__1841\ : IoSpan4Mux
    port map (
            O => \N__15416\,
            I => \N__15396\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__15413\,
            I => \N__15396\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__15410\,
            I => \N__15396\
        );

    \I__1838\ : IoInMux
    port map (
            O => \N__15409\,
            I => \N__15393\
        );

    \I__1837\ : IoInMux
    port map (
            O => \N__15408\,
            I => \N__15390\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15405\,
            I => \N__15387\
        );

    \I__1835\ : IoInMux
    port map (
            O => \N__15404\,
            I => \N__15384\
        );

    \I__1834\ : IoInMux
    port map (
            O => \N__15403\,
            I => \N__15381\
        );

    \I__1833\ : IoSpan4Mux
    port map (
            O => \N__15396\,
            I => \N__15374\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__15393\,
            I => \N__15374\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15374\
        );

    \I__1830\ : IoSpan4Mux
    port map (
            O => \N__15387\,
            I => \N__15365\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__15384\,
            I => \N__15365\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15365\
        );

    \I__1827\ : IoSpan4Mux
    port map (
            O => \N__15374\,
            I => \N__15359\
        );

    \I__1826\ : IoInMux
    port map (
            O => \N__15373\,
            I => \N__15356\
        );

    \I__1825\ : IoInMux
    port map (
            O => \N__15372\,
            I => \N__15353\
        );

    \I__1824\ : IoSpan4Mux
    port map (
            O => \N__15365\,
            I => \N__15349\
        );

    \I__1823\ : IoInMux
    port map (
            O => \N__15364\,
            I => \N__15346\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__15363\,
            I => \N__15343\
        );

    \I__1821\ : IoInMux
    port map (
            O => \N__15362\,
            I => \N__15340\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__15359\,
            I => \N__15337\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15334\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__15353\,
            I => \N__15331\
        );

    \I__1817\ : IoInMux
    port map (
            O => \N__15352\,
            I => \N__15328\
        );

    \I__1816\ : IoSpan4Mux
    port map (
            O => \N__15349\,
            I => \N__15323\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__15346\,
            I => \N__15323\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__15343\,
            I => \N__15320\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__15340\,
            I => \N__15317\
        );

    \I__1812\ : IoSpan4Mux
    port map (
            O => \N__15337\,
            I => \N__15312\
        );

    \I__1811\ : IoSpan4Mux
    port map (
            O => \N__15334\,
            I => \N__15312\
        );

    \I__1810\ : Span4Mux_s1_v
    port map (
            O => \N__15331\,
            I => \N__15308\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__15328\,
            I => \N__15305\
        );

    \I__1808\ : Span4Mux_s2_v
    port map (
            O => \N__15323\,
            I => \N__15302\
        );

    \I__1807\ : Span4Mux_s2_v
    port map (
            O => \N__15320\,
            I => \N__15299\
        );

    \I__1806\ : Span12Mux_s2_v
    port map (
            O => \N__15317\,
            I => \N__15296\
        );

    \I__1805\ : Span4Mux_s2_h
    port map (
            O => \N__15312\,
            I => \N__15293\
        );

    \I__1804\ : IoInMux
    port map (
            O => \N__15311\,
            I => \N__15290\
        );

    \I__1803\ : Sp12to4
    port map (
            O => \N__15308\,
            I => \N__15287\
        );

    \I__1802\ : IoSpan4Mux
    port map (
            O => \N__15305\,
            I => \N__15284\
        );

    \I__1801\ : Sp12to4
    port map (
            O => \N__15302\,
            I => \N__15279\
        );

    \I__1800\ : Sp12to4
    port map (
            O => \N__15299\,
            I => \N__15279\
        );

    \I__1799\ : Span12Mux_v
    port map (
            O => \N__15296\,
            I => \N__15276\
        );

    \I__1798\ : Sp12to4
    port map (
            O => \N__15293\,
            I => \N__15271\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__15290\,
            I => \N__15271\
        );

    \I__1796\ : Span12Mux_h
    port map (
            O => \N__15287\,
            I => \N__15268\
        );

    \I__1795\ : Span4Mux_s2_h
    port map (
            O => \N__15284\,
            I => \N__15265\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__15279\,
            I => \N__15262\
        );

    \I__1793\ : Span12Mux_v
    port map (
            O => \N__15276\,
            I => \N__15257\
        );

    \I__1792\ : Span12Mux_s10_h
    port map (
            O => \N__15271\,
            I => \N__15257\
        );

    \I__1791\ : Span12Mux_v
    port map (
            O => \N__15268\,
            I => \N__15252\
        );

    \I__1790\ : Sp12to4
    port map (
            O => \N__15265\,
            I => \N__15252\
        );

    \I__1789\ : Span12Mux_v
    port map (
            O => \N__15262\,
            I => \N__15247\
        );

    \I__1788\ : Span12Mux_h
    port map (
            O => \N__15257\,
            I => \N__15247\
        );

    \I__1787\ : Span12Mux_v
    port map (
            O => \N__15252\,
            I => \N__15244\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__15247\,
            I => dma_0_i
        );

    \I__1785\ : Odrv12
    port map (
            O => \N__15244\,
            I => dma_0_i
        );

    \I__1784\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__15227\,
            I => \this_ppu.oam_cache.mem_7\
        );

    \I__1779\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__15221\,
            I => \N__15218\
        );

    \I__1777\ : Span12Mux_h
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__15215\,
            I => \this_ppu.oam_cache.mem_3\
        );

    \I__1775\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__15209\,
            I => \M_this_oam_ram_write_data_5\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__15200\,
            I => \M_this_oam_ram_write_data_7\
        );

    \I__1770\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__15194\,
            I => \M_this_oam_ram_read_data_28\
        );

    \I__1768\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__1766\ : Span4Mux_v
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__15182\,
            I => \N__15179\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__15179\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_28\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__15173\,
            I => \M_this_oam_ram_read_data_29\
        );

    \I__1761\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__1759\ : Sp12to4
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__15161\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_29\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15158\,
            I => \N__15155\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__15155\,
            I => \N__15152\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__15152\,
            I => \M_this_oam_ram_write_data_16\
        );

    \I__1754\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15146\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__15146\,
            I => \N__15143\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__15143\,
            I => \M_this_oam_ram_write_data_22\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15137\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__1749\ : Span12Mux_s8_h
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__15131\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_19\
        );

    \I__1747\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15122\
        );

    \I__1746\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15122\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__15119\,
            I => \M_this_oam_ram_read_data_19\
        );

    \I__1743\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__15107\,
            I => \N__15104\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__15104\,
            I => \M_this_oam_ram_read_data_i_19\
        );

    \I__1738\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15098\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__15098\,
            I => \N__15095\
        );

    \I__1736\ : Span4Mux_v
    port map (
            O => \N__15095\,
            I => \N__15092\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__15092\,
            I => \N__15089\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__15089\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_20\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15083\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15083\,
            I => \M_this_oam_ram_write_data_13\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__15077\,
            I => \M_this_oam_ram_write_data_15\
        );

    \I__1729\ : InMux
    port map (
            O => \N__15074\,
            I => \N__15071\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15071\,
            I => \N__15068\
        );

    \I__1727\ : Span4Mux_s1_v
    port map (
            O => \N__15068\,
            I => \N__15065\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__15065\,
            I => \M_this_oam_ram_write_data_18\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15059\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__15059\,
            I => \N__15056\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__15056\,
            I => \M_this_oam_ram_read_data_31\
        );

    \I__1722\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__1720\ : Span4Mux_h
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__15041\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_31\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15038\,
            I => \N__15035\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__15035\,
            I => \M_this_oam_ram_write_data_8\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__15026\,
            I => \M_this_data_tmp_qZ0Z_3\
        );

    \I__1712\ : InMux
    port map (
            O => \N__15023\,
            I => \N__15020\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__15020\,
            I => \M_this_oam_ram_write_data_3\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__15010\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15007\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__15010\,
            I => \N__15004\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__15007\,
            I => \N__15001\
        );

    \I__1705\ : Odrv12
    port map (
            O => \N__15004\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__15001\,
            I => \M_this_oam_ram_read_data_21\
        );

    \I__1703\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14993\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__14990\,
            I => \M_this_oam_ram_read_data_i_21\
        );

    \I__1700\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14984\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14981\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__14981\,
            I => \M_this_data_tmp_qZ0Z_6\
        );

    \I__1697\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__14975\,
            I => \M_this_oam_ram_write_data_6\
        );

    \I__1695\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14966\
        );

    \I__1694\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14966\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14963\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__14963\,
            I => \N__14960\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__14957\,
            I => \M_this_oam_ram_read_data_22\
        );

    \I__1689\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__14951\,
            I => \M_this_oam_ram_read_data_i_22\
        );

    \I__1687\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14944\
        );

    \I__1686\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14941\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__14944\,
            I => \N__14936\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__14941\,
            I => \N__14936\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__14936\,
            I => \N__14933\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__14930\,
            I => \M_this_oam_ram_read_data_23\
        );

    \I__1680\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__14921\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_23\
        );

    \I__1677\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__1675\ : Span4Mux_v
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__14909\,
            I => \N__14906\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__14906\,
            I => \M_this_oam_ram_read_data_24\
        );

    \I__1672\ : InMux
    port map (
            O => \N__14903\,
            I => \N__14900\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__14897\,
            I => \N__14894\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__14894\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_24\
        );

    \I__1668\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__14882\,
            I => \N__14879\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__14879\,
            I => \M_this_oam_ram_read_data_25\
        );

    \I__1663\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__14873\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_25\
        );

    \I__1661\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__14867\,
            I => \N__14864\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__14858\,
            I => \M_this_oam_ram_read_data_26\
        );

    \I__1656\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__14849\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_26\
        );

    \I__1653\ : InMux
    port map (
            O => \N__14846\,
            I => \N__14843\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__14843\,
            I => \M_this_oam_ram_write_data_14\
        );

    \I__1651\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14837\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__14837\,
            I => \N__14834\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__14834\,
            I => \M_this_oam_ram_read_data_30\
        );

    \I__1648\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__1645\ : Span4Mux_v
    port map (
            O => \N__14822\,
            I => \N__14819\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__14819\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_30\
        );

    \I__1643\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__14813\,
            I => \this_ppu.M_this_oam_ram_read_data_i_17\
        );

    \I__1641\ : InMux
    port map (
            O => \N__14810\,
            I => \N__14807\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__14807\,
            I => \this_ppu.M_this_oam_ram_read_data_i_18\
        );

    \I__1639\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__14801\,
            I => \this_ppu.m28_e_i_o2_0\
        );

    \I__1637\ : InMux
    port map (
            O => \N__14798\,
            I => \this_ppu.un1_oam_data_1_cry_2\
        );

    \I__1636\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14792\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__14792\,
            I => \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\
        );

    \I__1634\ : InMux
    port map (
            O => \N__14789\,
            I => \this_ppu.un1_oam_data_1_cry_3\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__1632\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14780\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__14780\,
            I => \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\
        );

    \I__1630\ : InMux
    port map (
            O => \N__14777\,
            I => \this_ppu.un1_oam_data_1_cry_4\
        );

    \I__1629\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__14771\,
            I => \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\
        );

    \I__1627\ : InMux
    port map (
            O => \N__14768\,
            I => \this_ppu.un1_oam_data_1_cry_5\
        );

    \I__1626\ : InMux
    port map (
            O => \N__14765\,
            I => \this_ppu.un1_oam_data_1_cry_6\
        );

    \I__1625\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__14759\,
            I => \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0\
        );

    \I__1623\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__14753\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_21\
        );

    \I__1621\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__14747\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_22\
        );

    \I__1619\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__14738\,
            I => \this_ppu.oam_cache.mem_18\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__1615\ : CascadeBuf
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__1613\ : InMux
    port map (
            O => \N__14726\,
            I => \N__14723\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__14723\,
            I => \this_ppu.N_777_0\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__1610\ : CascadeBuf
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__1608\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14708\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__14708\,
            I => \this_ppu.N_776_0\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__14705\,
            I => \this_ppu.N_932_0_cascade_\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \this_ppu.un1_M_state_q_7_i_0_0_cascade_\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__1603\ : CascadeBuf
    port map (
            O => \N__14696\,
            I => \N__14693\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__1601\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__14687\,
            I => \this_ppu.N_775_0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__14681\,
            I => \this_ppu.N_932_0\
        );

    \I__1597\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14672\
        );

    \I__1596\ : InMux
    port map (
            O => \N__14677\,
            I => \N__14672\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__1594\ : Span12Mux_v
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__1593\ : Odrv12
    port map (
            O => \N__14666\,
            I => \this_ppu.N_838_7\
        );

    \I__1592\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__14660\,
            I => \this_ppu.M_this_oam_ram_read_data_i_16\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \this_vga_ramdac.m16_cascade_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__14645\,
            I => \N__14641\
        );

    \I__1585\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14638\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__14641\,
            I => \this_vga_ramdac.N_3141_reto\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__14638\,
            I => \this_vga_ramdac.N_3141_reto\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \this_vga_ramdac.m19_cascade_\
        );

    \I__1581\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__14621\,
            I => \N__14617\
        );

    \I__1577\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__14617\,
            I => \this_vga_ramdac.N_3142_reto\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__14614\,
            I => \this_vga_ramdac.N_3142_reto\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14599\
        );

    \I__1573\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14599\
        );

    \I__1572\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14590\
        );

    \I__1571\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14590\
        );

    \I__1570\ : InMux
    port map (
            O => \N__14605\,
            I => \N__14590\
        );

    \I__1569\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14590\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__14599\,
            I => \M_this_vram_read_data_0\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__14590\,
            I => \M_this_vram_read_data_0\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__1565\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14575\
        );

    \I__1564\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14566\
        );

    \I__1563\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14566\
        );

    \I__1562\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14566\
        );

    \I__1561\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14566\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__14575\,
            I => \M_this_vram_read_data_2\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__14566\,
            I => \M_this_vram_read_data_2\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \N__14553\
        );

    \I__1557\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14548\
        );

    \I__1556\ : InMux
    port map (
            O => \N__14559\,
            I => \N__14548\
        );

    \I__1555\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14539\
        );

    \I__1554\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14539\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14539\
        );

    \I__1552\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14539\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__14548\,
            I => \M_this_vram_read_data_3\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__14539\,
            I => \M_this_vram_read_data_3\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__14534\,
            I => \N__14527\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__14533\,
            I => \N__14524\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__14532\,
            I => \N__14521\
        );

    \I__1546\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14515\
        );

    \I__1545\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14515\
        );

    \I__1544\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14506\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14506\
        );

    \I__1542\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14506\
        );

    \I__1541\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14506\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__14515\,
            I => \M_this_vram_read_data_1\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__14506\,
            I => \M_this_vram_read_data_1\
        );

    \I__1538\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14498\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__14495\,
            I => \N__14492\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__14492\,
            I => \this_vga_ramdac.m6\
        );

    \I__1534\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__14483\,
            I => \N__14480\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__14480\,
            I => \this_ppu.oam_cache.mem_17\
        );

    \I__1530\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14474\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__14474\,
            I => \this_ppu.oam_cache.M_oam_cache_read_data_17\
        );

    \I__1528\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__14468\,
            I => \N__14465\
        );

    \I__1526\ : Span4Mux_v
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__14462\,
            I => \this_ppu.oam_cache.mem_16\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__14456\,
            I => \this_vga_ramdac.i2_mux_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14450\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14447\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__14447\,
            I => \N__14443\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__14446\,
            I => \N__14440\
        );

    \I__1518\ : Span4Mux_h
    port map (
            O => \N__14443\,
            I => \N__14437\
        );

    \I__1517\ : InMux
    port map (
            O => \N__14440\,
            I => \N__14434\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__14437\,
            I => \this_vga_ramdac.N_3143_reto\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__14434\,
            I => \this_vga_ramdac.N_3143_reto\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__14429\,
            I => \this_vga_ramdac.i2_mux_cascade_\
        );

    \I__1513\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14419\
        );

    \I__1511\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14416\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__14419\,
            I => \N__14411\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14411\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__14411\,
            I => \this_vga_ramdac.N_3140_reto\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__14408\,
            I => \this_vga_ramdac.N_24_mux_cascade_\
        );

    \I__1506\ : InMux
    port map (
            O => \N__14405\,
            I => \N__14402\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__14399\,
            I => \N__14395\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14392\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__14395\,
            I => \this_vga_ramdac.N_3138_reto\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__14392\,
            I => \this_vga_ramdac.N_3138_reto\
        );

    \I__1500\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14384\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14381\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__14378\,
            I => \this_ppu.oam_cache.mem_6\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__14375\,
            I => \N__14371\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14365\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14365\
        );

    \I__1493\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14362\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14365\,
            I => \N__14355\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14352\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__14361\,
            I => \N__14346\
        );

    \I__1489\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14342\
        );

    \I__1488\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14339\
        );

    \I__1487\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14336\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__14355\,
            I => \N__14331\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__14352\,
            I => \N__14331\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14326\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14326\
        );

    \I__1482\ : InMux
    port map (
            O => \N__14349\,
            I => \N__14319\
        );

    \I__1481\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14319\
        );

    \I__1480\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14319\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__14342\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14339\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14336\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__14331\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__14326\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__14319\,
            I => \this_vga_signals.M_hcounter_qZ0Z_5\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \N__14303\
        );

    \I__1472\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14300\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__14300\,
            I => \this_vga_signals.M_hcounter_d7lt7_0\
        );

    \I__1470\ : InMux
    port map (
            O => \N__14297\,
            I => \N__14287\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14296\,
            I => \N__14287\
        );

    \I__1468\ : InMux
    port map (
            O => \N__14295\,
            I => \N__14287\
        );

    \I__1467\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14284\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__14287\,
            I => \N__14280\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14277\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14269\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__14280\,
            I => \N__14264\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__14277\,
            I => \N__14264\
        );

    \I__1461\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14257\
        );

    \I__1460\ : InMux
    port map (
            O => \N__14275\,
            I => \N__14257\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14257\
        );

    \I__1458\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14252\
        );

    \I__1457\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14252\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__14269\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__14264\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__14257\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__14252\,
            I => \this_vga_signals.M_hcounter_qZ0Z_6\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__14243\,
            I => \N__14237\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14234\
        );

    \I__1450\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14231\
        );

    \I__1449\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14226\
        );

    \I__1448\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14226\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14221\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__14231\,
            I => \N__14221\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__14226\,
            I => \N__14213\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__14221\,
            I => \N__14210\
        );

    \I__1443\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14205\
        );

    \I__1442\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14205\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \N__14202\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__14217\,
            I => \N__14199\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14196\
        );

    \I__1438\ : Span4Mux_h
    port map (
            O => \N__14213\,
            I => \N__14189\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__14210\,
            I => \N__14189\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14205\,
            I => \N__14189\
        );

    \I__1435\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14186\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14183\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__14196\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1432\ : Odrv4
    port map (
            O => \N__14189\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__14186\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__14183\,
            I => \this_vga_signals.M_hcounter_qZ0Z_9\
        );

    \I__1429\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14166\
        );

    \I__1428\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14166\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14162\
        );

    \I__1426\ : InMux
    port map (
            O => \N__14171\,
            I => \N__14159\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__14166\,
            I => \N__14156\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14153\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__14162\,
            I => \N__14150\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__14159\,
            I => \N__14146\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__14156\,
            I => \N__14141\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__14153\,
            I => \N__14141\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__14150\,
            I => \N__14136\
        );

    \I__1418\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14133\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__14146\,
            I => \N__14130\
        );

    \I__1416\ : Span4Mux_h
    port map (
            O => \N__14141\,
            I => \N__14127\
        );

    \I__1415\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14124\
        );

    \I__1414\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14121\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__14136\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__14133\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1411\ : Odrv4
    port map (
            O => \N__14130\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__14127\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__14124\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__14121\,
            I => \this_vga_signals.M_hcounter_qZ0Z_8\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__14108\,
            I => \this_vga_signals.N_864_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14105\,
            I => \N__14094\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14094\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14094\
        );

    \I__1403\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14090\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14087\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__14094\,
            I => \N__14084\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14081\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__14090\,
            I => \N__14078\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__14087\,
            I => \N__14074\
        );

    \I__1397\ : Span4Mux_h
    port map (
            O => \N__14084\,
            I => \N__14069\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__14081\,
            I => \N__14069\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__14078\,
            I => \N__14064\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14061\
        );

    \I__1393\ : Span4Mux_h
    port map (
            O => \N__14074\,
            I => \N__14058\
        );

    \I__1392\ : Span4Mux_h
    port map (
            O => \N__14069\,
            I => \N__14055\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14052\
        );

    \I__1390\ : InMux
    port map (
            O => \N__14067\,
            I => \N__14049\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__14064\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__14061\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__14058\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__14055\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14052\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__14049\,
            I => \this_vga_signals.M_hcounter_qZ0Z_7\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14033\,
            I => \N__14029\
        );

    \I__1381\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__1380\ : Span4Mux_v
    port map (
            O => \N__14029\,
            I => \N__14021\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__14026\,
            I => \N__14021\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__14021\,
            I => \M_this_oam_ram_read_data_5\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14015\,
            I => \N__14011\
        );

    \I__1375\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__14011\,
            I => \N__14003\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__14008\,
            I => \N__14003\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__14003\,
            I => \M_this_oam_ram_read_data_2\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__14000\,
            I => \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__13994\,
            I => \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4\
        );

    \I__1368\ : CascadeMux
    port map (
            O => \N__13991\,
            I => \this_ppu.m35_i_a2_3_cascade_\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \this_ppu.N_802_cascade_\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__13985\,
            I => \N__13980\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13977\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__13983\,
            I => \N__13974\
        );

    \I__1363\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13969\
        );

    \I__1362\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13961\
        );

    \I__1361\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13961\
        );

    \I__1360\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13961\
        );

    \I__1359\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13956\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__13969\,
            I => \N__13953\
        );

    \I__1357\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13950\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__13961\,
            I => \N__13947\
        );

    \I__1355\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13944\
        );

    \I__1354\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13941\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13930\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__13953\,
            I => \N__13930\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__13950\,
            I => \N__13930\
        );

    \I__1350\ : Span4Mux_v
    port map (
            O => \N__13947\,
            I => \N__13930\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__13944\,
            I => \N__13930\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__13941\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__13930\,
            I => \this_vga_signals.M_hcounter_qZ0Z_3\
        );

    \I__1346\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13921\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__13924\,
            I => \N__13918\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__13921\,
            I => \N__13912\
        );

    \I__1343\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13906\
        );

    \I__1342\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13906\
        );

    \I__1341\ : InMux
    port map (
            O => \N__13916\,
            I => \N__13901\
        );

    \I__1340\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13901\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__13912\,
            I => \N__13896\
        );

    \I__1338\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13893\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__13906\,
            I => \N__13888\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__13901\,
            I => \N__13888\
        );

    \I__1335\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13885\
        );

    \I__1334\ : InMux
    port map (
            O => \N__13899\,
            I => \N__13882\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__13896\,
            I => \N__13873\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__13893\,
            I => \N__13873\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__13888\,
            I => \N__13873\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__13885\,
            I => \N__13873\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__13882\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__13873\,
            I => \this_vga_signals.M_hcounter_qZ0Z_2\
        );

    \I__1327\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__13865\,
            I => \N__13862\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__1324\ : Span4Mux_h
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__13856\,
            I => \this_vga_signals.un2_hsynclto3_1\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__13853\,
            I => \this_vga_signals.un2_hsynclto3_1_cascade_\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \N__13847\
        );

    \I__1320\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13841\
        );

    \I__1319\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13835\
        );

    \I__1318\ : InMux
    port map (
            O => \N__13845\,
            I => \N__13835\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__13844\,
            I => \N__13832\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__13841\,
            I => \N__13827\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__13840\,
            I => \N__13822\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__13835\,
            I => \N__13818\
        );

    \I__1313\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13813\
        );

    \I__1312\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13813\
        );

    \I__1311\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13810\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__13827\,
            I => \N__13807\
        );

    \I__1309\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13804\
        );

    \I__1308\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13797\
        );

    \I__1307\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13797\
        );

    \I__1306\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13797\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__13818\,
            I => \N__13790\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__13813\,
            I => \N__13790\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__13810\,
            I => \N__13790\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__13807\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__13804\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__13797\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__13790\,
            I => \this_vga_signals.M_hcounter_qZ0Z_4\
        );

    \I__1298\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13778\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__13778\,
            I => \N__13772\
        );

    \I__1296\ : InMux
    port map (
            O => \N__13777\,
            I => \N__13769\
        );

    \I__1295\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13764\
        );

    \I__1294\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13761\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__13772\,
            I => \N__13755\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__13769\,
            I => \N__13755\
        );

    \I__1291\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13752\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__13767\,
            I => \N__13749\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__13764\,
            I => \N__13744\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13744\
        );

    \I__1287\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13741\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__13755\,
            I => \N__13736\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13736\
        );

    \I__1284\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13733\
        );

    \I__1283\ : Span12Mux_v
    port map (
            O => \N__13744\,
            I => \N__13728\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13728\
        );

    \I__1281\ : Span4Mux_h
    port map (
            O => \N__13736\,
            I => \N__13725\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13722\
        );

    \I__1279\ : Odrv12
    port map (
            O => \N__13728\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__13725\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__13722\,
            I => \this_vga_ramdac.M_this_vga_ramdac_en_reto\
        );

    \I__1276\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13712\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__13712\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__1273\ : CascadeBuf
    port map (
            O => \N__13706\,
            I => \N__13701\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__13705\,
            I => \N__13697\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__13704\,
            I => \N__13694\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__13701\,
            I => \N__13691\
        );

    \I__1269\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13688\
        );

    \I__1268\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13683\
        );

    \I__1267\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13683\
        );

    \I__1266\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13680\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__13688\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_3\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__13683\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_3\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__13680\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_3\
        );

    \I__1262\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__13670\,
            I => \this_ppu.oam_cache.N_826_0\
        );

    \I__1260\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13661\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__13658\,
            I => \this_ppu.oam_cache.N_824_0\
        );

    \I__1256\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__1254\ : Span4Mux_h
    port map (
            O => \N__13649\,
            I => \N__13646\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__13646\,
            I => \this_ppu.oam_cache.N_821_0\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__1250\ : Span4Mux_h
    port map (
            O => \N__13637\,
            I => \N__13634\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__13634\,
            I => \this_ppu.oam_cache.N_822_0\
        );

    \I__1248\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13628\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__13628\,
            I => \N__13625\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__13622\,
            I => \this_ppu.oam_cache.N_819_0\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13616\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__1242\ : Span4Mux_h
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__13610\,
            I => \N__13607\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__13607\,
            I => \this_ppu.oam_cache.N_825_0\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__13601\,
            I => \N__13598\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__13598\,
            I => \N__13594\
        );

    \I__1236\ : InMux
    port map (
            O => \N__13597\,
            I => \N__13591\
        );

    \I__1235\ : Span4Mux_v
    port map (
            O => \N__13594\,
            I => \N__13586\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__13591\,
            I => \N__13586\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__13586\,
            I => \M_this_oam_ram_read_data_0\
        );

    \I__1232\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13576\
        );

    \I__1230\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13573\
        );

    \I__1229\ : Span12Mux_s7_h
    port map (
            O => \N__13576\,
            I => \N__13570\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__13573\,
            I => \N__13567\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__13570\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__13567\,
            I => \M_this_oam_ram_read_data_6\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13562\,
            I => \N__13558\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__13561\,
            I => \N__13555\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13552\
        );

    \I__1222\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13549\
        );

    \I__1221\ : Span4Mux_v
    port map (
            O => \N__13552\,
            I => \N__13544\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13544\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__13544\,
            I => \M_this_oam_ram_read_data_1\
        );

    \I__1218\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__13538\,
            I => \N__13535\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__13535\,
            I => \N__13531\
        );

    \I__1215\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13528\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__13531\,
            I => \N__13523\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__13528\,
            I => \N__13523\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__13523\,
            I => \M_this_oam_ram_read_data_3\
        );

    \I__1211\ : InMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__13517\,
            I => \N__13513\
        );

    \I__1209\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13510\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__13513\,
            I => \N__13505\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13505\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__13505\,
            I => \M_this_oam_ram_read_data_7\
        );

    \I__1205\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13499\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__13499\,
            I => \N__13495\
        );

    \I__1203\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13492\
        );

    \I__1202\ : Span4Mux_v
    port map (
            O => \N__13495\,
            I => \N__13487\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__13492\,
            I => \N__13487\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__13487\,
            I => \M_this_oam_ram_read_data_4\
        );

    \I__1199\ : InMux
    port map (
            O => \N__13484\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\
        );

    \I__1198\ : InMux
    port map (
            O => \N__13481\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\
        );

    \I__1197\ : InMux
    port map (
            O => \N__13478\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_3\
        );

    \I__1196\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13471\
        );

    \I__1195\ : InMux
    port map (
            O => \N__13474\,
            I => \N__13468\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__13471\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_4\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__13468\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_4\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__13463\,
            I => \this_ppu.m71_i_o2_0_cascade_\
        );

    \I__1191\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__13457\,
            I => \this_ppu.m71_i_o2_1\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \N__13451\
        );

    \I__1188\ : CascadeBuf
    port map (
            O => \N__13451\,
            I => \N__13446\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__13450\,
            I => \N__13443\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__13449\,
            I => \N__13439\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__13446\,
            I => \N__13436\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13443\,
            I => \N__13431\
        );

    \I__1183\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13431\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13428\
        );

    \I__1181\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13425\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__13431\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_0\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__13428\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_0\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__13425\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_0\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__13415\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__1174\ : CascadeBuf
    port map (
            O => \N__13409\,
            I => \N__13404\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__13408\,
            I => \N__13401\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__13407\,
            I => \N__13397\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__13404\,
            I => \N__13394\
        );

    \I__1170\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13391\
        );

    \I__1169\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13386\
        );

    \I__1168\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13386\
        );

    \I__1167\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13383\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__13391\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__13386\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__13383\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_2\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__1162\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13370\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__13370\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__1159\ : CascadeBuf
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__13361\,
            I => \N__13355\
        );

    \I__1157\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13352\
        );

    \I__1156\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13349\
        );

    \I__1155\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13346\
        );

    \I__1154\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13343\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__13352\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__13349\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__13346\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__13343\,
            I => \this_ppu.M_oam_cache_cnt_qZ0Z_1\
        );

    \I__1149\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13331\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__13325\,
            I => \N__13322\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__13322\,
            I => \M_this_oam_ram_read_data_14\
        );

    \I__1144\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13316\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__13316\,
            I => \N__13313\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__13313\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_14\
        );

    \I__1141\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__13307\,
            I => \N__13304\
        );

    \I__1139\ : Span4Mux_v
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__13301\,
            I => \N__13298\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__13298\,
            I => \M_this_oam_ram_read_data_15\
        );

    \I__1136\ : InMux
    port map (
            O => \N__13295\,
            I => \N__13292\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__13292\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_15\
        );

    \I__1134\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__13286\,
            I => \this_ppu.oam_cache.N_823_0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__13280\,
            I => \this_ppu.oam_cache.N_820_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__1126\ : Span4Mux_v
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__13262\,
            I => \M_this_oam_ram_read_data_8\
        );

    \I__1124\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__13256\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_8\
        );

    \I__1122\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__13247\,
            I => \N__13244\
        );

    \I__1119\ : Sp12to4
    port map (
            O => \N__13244\,
            I => \N__13241\
        );

    \I__1118\ : Odrv12
    port map (
            O => \N__13241\,
            I => \M_this_oam_ram_read_data_9\
        );

    \I__1117\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__13235\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_9\
        );

    \I__1115\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__1113\ : Span12Mux_v
    port map (
            O => \N__13226\,
            I => \N__13223\
        );

    \I__1112\ : Odrv12
    port map (
            O => \N__13223\,
            I => \M_this_oam_ram_read_data_10\
        );

    \I__1111\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__13217\,
            I => \this_ppu.oam_cache.M_oam_cache_write_data_10\
        );

    \I__1109\ : InMux
    port map (
            O => \N__13214\,
            I => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\
        );

    \I__1108\ : InMux
    port map (
            O => \N__13211\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_1\
        );

    \I__1107\ : InMux
    port map (
            O => \N__13208\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_2\
        );

    \I__1106\ : InMux
    port map (
            O => \N__13205\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_3\
        );

    \I__1105\ : InMux
    port map (
            O => \N__13202\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_4\
        );

    \I__1104\ : InMux
    port map (
            O => \N__13199\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_5\
        );

    \I__1103\ : InMux
    port map (
            O => \N__13196\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_6\
        );

    \I__1102\ : InMux
    port map (
            O => \N__13193\,
            I => \this_vga_signals.un1_M_hcounter_d_cry_7\
        );

    \I__1101\ : InMux
    port map (
            O => \N__13190\,
            I => \bfn_7_18_0_\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\
        );

    \I__1099\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13180\
        );

    \I__1098\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13177\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__13180\,
            I => \this_vga_signals.mult1_un68_sum_c3_2\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__13177\,
            I => \this_vga_signals.mult1_un68_sum_c3_2\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__13172\,
            I => \this_vga_signals.mult1_un68_sum_c3_2_cascade_\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__1093\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13163\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__13163\,
            I => \N__13160\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__13160\,
            I => \N__13157\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__13157\,
            I => \M_this_vga_signals_address_3\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__1088\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__13142\,
            I => \M_this_vga_signals_address_5\
        );

    \I__1084\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13135\
        );

    \I__1083\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13132\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__13135\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__13132\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__1079\ : InMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__13121\,
            I => \N__13118\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__13118\,
            I => \N__13115\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__13115\,
            I => \M_this_vga_signals_address_4\
        );

    \I__1075\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13106\
        );

    \I__1074\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13099\
        );

    \I__1073\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13099\
        );

    \I__1072\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13099\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__13106\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__13099\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__13094\,
            I => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\
        );

    \I__1068\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13087\
        );

    \I__1067\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13084\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__13087\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__13084\,
            I => \this_vga_signals.SUM_3\
        );

    \I__1064\ : InMux
    port map (
            O => \N__13079\,
            I => \N__13076\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__13076\,
            I => \this_vga_signals.mult1_un54_sum_c3_0\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\
        );

    \I__1061\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13067\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__13067\,
            I => \this_vga_signals.if_m1_1\
        );

    \I__1059\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13057\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__13060\,
            I => \N__13054\
        );

    \I__1056\ : Span4Mux_h
    port map (
            O => \N__13057\,
            I => \N__13051\
        );

    \I__1055\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13048\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__13051\,
            I => \this_vga_ramdac.N_3139_reto\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__13048\,
            I => \this_vga_ramdac.N_3139_reto\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__13043\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\
        );

    \I__1051\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13030\
        );

    \I__1050\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13030\
        );

    \I__1049\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13030\
        );

    \I__1048\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13027\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__13030\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__13027\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__13022\,
            I => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__13019\,
            I => \N__13016\
        );

    \I__1043\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13013\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__13013\,
            I => \N__13010\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__13010\,
            I => \M_this_vga_signals_address_2\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__13007\,
            I => \this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_\
        );

    \I__1039\ : InMux
    port map (
            O => \N__13004\,
            I => \N__13001\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__13001\,
            I => \this_vga_signals.if_m7_0_o4_1_ns_1\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__12998\,
            I => \this_vga_signals.SUM_3_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__12992\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_1\
        );

    \I__1034\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12986\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__12986\,
            I => \this_vga_signals.mult1_un89_sum_c3_0\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__1031\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12977\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__12974\,
            I => \M_this_vga_signals_address_0\
        );

    \I__1028\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12967\
        );

    \I__1027\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__12967\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__12964\,
            I => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\
        );

    \I__1024\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12956\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__12956\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1_2\
        );

    \I__1022\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__12950\,
            I => \this_vga_signals.un2_hsynclto6_0\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__12947\,
            I => \this_vga_signals.un4_hsynclt7_cascade_\
        );

    \I__1019\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12941\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__12941\,
            I => \this_vga_signals.hsync_1_1\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__12938\,
            I => \this_vga_signals.un4_hsynclt8_0_cascade_\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__12935\,
            I => \N__12932\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__1014\ : Span12Mux_s2_v
    port map (
            O => \N__12929\,
            I => \N__12926\
        );

    \I__1013\ : Span12Mux_v
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__1012\ : Odrv12
    port map (
            O => \N__12923\,
            I => this_vga_signals_hsync_1_i
        );

    \I__1011\ : IoInMux
    port map (
            O => \N__12920\,
            I => \N__12917\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__12917\,
            I => \N__12914\
        );

    \I__1009\ : Span4Mux_s0_v
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__1007\ : Span4Mux_v
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__1006\ : Span4Mux_v
    port map (
            O => \N__12905\,
            I => \N__12902\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__12902\,
            I => this_vga_signals_hvisibility_i
        );

    \I__1004\ : IoInMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__12896\,
            I => \N__12893\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__12893\,
            I => this_vga_signals_vvisibility_i
        );

    \I__1001\ : IoInMux
    port map (
            O => \N__12890\,
            I => \N__12887\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__999\ : Span4Mux_s1_h
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__998\ : Sp12to4
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__997\ : Span12Mux_v
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__996\ : Odrv12
    port map (
            O => \N__12875\,
            I => rgb_c_0
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__12872\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_\
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__12869\,
            I => \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\
        );

    \I__993\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__12863\,
            I => \this_vga_signals.mult1_un89_sum_c3_1\
        );

    \I__991\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12854\
        );

    \I__990\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12854\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__12854\,
            I => \this_vga_signals.mult1_un82_sum_c3_0\
        );

    \I__988\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12845\
        );

    \I__987\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12845\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__12845\,
            I => \this_vga_signals.mult1_un82_sum_axbxc3_1\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__12842\,
            I => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__12839\,
            I => \N__12836\
        );

    \I__983\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12830\
        );

    \I__981\ : Odrv12
    port map (
            O => \N__12830\,
            I => \M_this_vga_signals_address_1\
        );

    \I__980\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__12824\,
            I => \this_vga_signals.SUM_3_1\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__977\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12812\
        );

    \I__976\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12812\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__12812\,
            I => \this_vga_signals.mult1_un75_sum_axb1\
        );

    \I__974\ : IoInMux
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12803\
        );

    \I__972\ : IoSpan4Mux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__971\ : IoSpan4Mux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__970\ : Span4Mux_s1_h
    port map (
            O => \N__12797\,
            I => \N__12794\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__12794\,
            I => rgb_c_3
        );

    \I__968\ : IoInMux
    port map (
            O => \N__12791\,
            I => \N__12788\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__12788\,
            I => \N__12785\
        );

    \I__966\ : Odrv12
    port map (
            O => \N__12785\,
            I => rgb_c_1
        );

    \I__965\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__12779\,
            I => \this_delay_clk.M_pipe_qZ0Z_1\
        );

    \I__963\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__12773\,
            I => \this_delay_clk.M_pipe_qZ0Z_2\
        );

    \I__961\ : IoInMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__959\ : Odrv12
    port map (
            O => \N__12764\,
            I => rgb_c_2
        );

    \I__958\ : IoInMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__956\ : Span4Mux_s3_h
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__955\ : Span4Mux_v
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__12746\,
            I => rgb_c_4
        );

    \I__952\ : IoInMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__12740\,
            I => \N__12737\
        );

    \I__950\ : Span4Mux_s3_h
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__12731\,
            I => rgb_c_5
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__946\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12722\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__12719\,
            I => \M_this_vga_signals_address_6\
        );

    \I__943\ : IoInMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__12713\,
            I => port_data_rw_0_i
        );

    \I__941\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__12707\,
            I => \N__12704\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__12704\,
            I => \N__12701\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__12701\,
            I => port_clk_c
        );

    \I__937\ : InMux
    port map (
            O => \N__12698\,
            I => \N__12695\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__12695\,
            I => \this_delay_clk.M_pipe_qZ0Z_0\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_ppu.un1_M_surface_y_d_cry_6\,
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_8\,
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_16\,
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_warmup_d_cry_24\,
            carryinitout => \bfn_10_23_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            carryinitout => \bfn_7_18_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_7_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_20_0_\
        );

    \IN_MUX_bfv_15_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_19_0_\
        );

    \IN_MUX_bfv_15_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \M_this_data_count_q_cry_7\,
            carryinitout => \bfn_15_20_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_21_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_24_0_\
        );

    \IN_MUX_bfv_21_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_ext_address_q_cry_7\,
            carryinitout => \bfn_21_25_0_\
        );

    \IN_MUX_bfv_9_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_21_0_\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_spr_address_q_cry_7\,
            carryinitout => \bfn_17_13_0_\
        );

    \IN_MUX_bfv_26_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_25_0_\
        );

    \IN_MUX_bfv_26_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \un1_M_this_map_address_q_cry_7\,
            carryinitout => \bfn_26_26_0_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNINK957_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__29654\,
            GLOBALBUFFEROUTPUT => \this_vga_signals.N_1188_g\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__31013\,
            GLOBALBUFFEROUTPUT => \M_this_reset_cond_out_g_0\
        );

    \this_reset_cond.M_stage_q_RNIC5C7_0_9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__30125\,
            GLOBALBUFFEROUTPUT => \N_527_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \this_vga_signals.port_data_rw_0_i_LC_1_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__34178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31540\,
            lcout => port_data_rw_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_1_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12698\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_0_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIQ1FH_3_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14654\,
            in2 => \_gnd_net_\,
            in3 => \N__13776\,
            lcout => rgb_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIOVEH_1_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13064\,
            lcout => rgb_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_3_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12776\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_2_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12782\,
            lcout => \this_delay_clk.M_pipe_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIP0FH_2_LC_4_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13760\,
            lcout => rgb_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_0_LC_4_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__15596\,
            in1 => \N__13868\,
            in2 => \N__13850\,
            in3 => \N__15539\,
            lcout => \this_vga_signals.un2_hsynclto6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIR2FH_4_LC_4_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14630\,
            lcout => rgb_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNIS3FH_5_LC_4_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14453\,
            lcout => rgb_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIFI285_9_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12827\,
            in2 => \_gnd_net_\,
            in3 => \N__26468\,
            lcout => \M_this_vga_signals_address_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__13917\,
            in1 => \N__13184\,
            in2 => \N__13985\,
            in3 => \N__12959\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1\,
            ltout => \this_vga_signals.mult1_un82_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_1_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001000010"
        )
    port map (
            in0 => \N__15581\,
            in1 => \N__15531\,
            in2 => \N__12872\,
            in3 => \N__12859\,
            lcout => \this_vga_signals.mult1_un89_sum_c3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_0_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001001001011"
        )
    port map (
            in0 => \N__13039\,
            in1 => \N__15582\,
            in2 => \N__12821\,
            in3 => \N__13916\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un89_sum_axbxc3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_axbxc3_1_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12850\,
            in2 => \N__12869\,
            in3 => \N__12860\,
            lcout => \this_vga_signals.mult1_un89_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un89_sum_c3_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010110"
        )
    port map (
            in0 => \N__13040\,
            in1 => \N__15583\,
            in2 => \N__13924\,
            in3 => \N__12866\,
            lcout => \this_vga_signals.mult1_un89_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_c3_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101110001001"
        )
    port map (
            in0 => \N__13915\,
            in1 => \N__12817\,
            in2 => \N__15591\,
            in3 => \N__13038\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un82_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNISNQ4B1_9_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__12851\,
            in1 => \_gnd_net_\,
            in2 => \N__12842\,
            in3 => \N__26469\,
            lcout => \M_this_vga_signals_address_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_9_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111010111"
        )
    port map (
            in0 => \N__14173\,
            in1 => \N__14103\,
            in2 => \N__14243\,
            in3 => \N__14295\,
            lcout => \this_vga_signals.SUM_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axb1_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13973\,
            in2 => \_gnd_net_\,
            in3 => \N__13183\,
            lcout => \this_vga_signals.mult1_un75_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un82_sum_axbxc3_1_2_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13845\,
            in1 => \N__13138\,
            in2 => \N__13983\,
            in3 => \N__13037\,
            lcout => \this_vga_signals.mult1_un82_sum_axbxc3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIKCQ82_7_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__12953\,
            in1 => \N__14104\,
            in2 => \N__14375\,
            in3 => \N__14296\,
            lcout => \this_vga_signals.hsync_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI62D41_1_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__13846\,
            in1 => \N__15592\,
            in2 => \N__13984\,
            in3 => \N__13925\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNIL6NV1_7_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14374\,
            in1 => \N__14105\,
            in2 => \N__12947\,
            in3 => \N__14297\,
            lcout => OPEN,
            ltout => \this_vga_signals.un4_hsynclt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI1FBO4_9_LC_5_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__12944\,
            in1 => \N__14240\,
            in2 => \N__12938\,
            in3 => \N__14174\,
            lcout => this_vga_signals_hsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNICT164_9_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__14241\,
            in1 => \N__14171\,
            in2 => \N__29618\,
            in3 => \N__14101\,
            lcout => \M_this_vga_ramdac_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIU8TO_9_LC_5_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__14102\,
            in1 => \N__14242\,
            in2 => \_gnd_net_\,
            in3 => \N__14172\,
            lcout => this_vga_signals_hvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_0_9_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29617\,
            lcout => this_vga_signals_vvisibility_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_RNINUEH_0_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14405\,
            lcout => rgb_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_1_LC_6_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011010110"
        )
    port map (
            in0 => \N__14359\,
            in1 => \N__12970\,
            in2 => \N__13844\,
            in3 => \N__13111\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un75_sum_axbxc3_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101000011010"
        )
    port map (
            in0 => \N__13968\,
            in1 => \N__13899\,
            in2 => \N__13043\,
            in3 => \N__13004\,
            lcout => \this_vga_signals.mult1_un75_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIUG6BC_9_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__26481\,
            in1 => \_gnd_net_\,
            in2 => \N__13022\,
            in3 => \_gnd_net_\,
            lcout => \M_this_vga_signals_address_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_1_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110101"
        )
    port map (
            in0 => \N__13110\,
            in1 => \_gnd_net_\,
            in2 => \N__14361\,
            in3 => \N__13831\,
            lcout => OPEN,
            ltout => \this_vga_signals.if_m7_0_o4_1_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m7_0_o4_1_ns_1_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010101011110"
        )
    port map (
            in0 => \N__14276\,
            in1 => \N__14349\,
            in2 => \N__13007\,
            in3 => \N__13091\,
            lcout => \this_vga_signals.if_m7_0_o4_1_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_0_9_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010111010111"
        )
    port map (
            in0 => \N__14140\,
            in1 => \N__14068\,
            in2 => \N__14218\,
            in3 => \N__14274\,
            lcout => \this_vga_signals.SUM_3\,
            ltout => \this_vga_signals.SUM_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_1_0_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011110"
        )
    port map (
            in0 => \N__14275\,
            in1 => \N__14345\,
            in2 => \N__12998\,
            in3 => \N__13109\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI73OIC3_9_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__12995\,
            in1 => \N__26480\,
            in2 => \_gnd_net_\,
            in3 => \N__12989\,
            lcout => \M_this_vga_signals_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un61_sum_axbxc3_2_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111000100110"
        )
    port map (
            in0 => \N__14358\,
            in1 => \N__12971\,
            in2 => \N__13840\,
            in3 => \N__13112\,
            lcout => \this_vga_signals.mult1_un61_sum_axbxc3_2\,
            ltout => \this_vga_signals.mult1_un61_sum_axbxc3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un68_sum_c3_0_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110101000000"
        )
    port map (
            in0 => \N__13959\,
            in1 => \N__13825\,
            in2 => \N__13187\,
            in3 => \N__13070\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_2\,
            ltout => \this_vga_signals.mult1_un68_sum_c3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI0J6BC_9_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13172\,
            in3 => \N__26460\,
            lcout => \M_this_vga_signals_address_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIRU9S6_9_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13079\,
            lcout => \M_this_vga_signals_address_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI59HG8_9_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26461\,
            in2 => \_gnd_net_\,
            in3 => \N__13139\,
            lcout => \M_this_vga_signals_address_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNI3L021_1_9_LC_6_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010111101"
        )
    port map (
            in0 => \N__14139\,
            in1 => \N__14067\,
            in2 => \N__14217\,
            in3 => \N__14272\,
            lcout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9\,
            ltout => \this_vga_signals.M_hcounter_q_esr_RNI3L021_1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_generate_plus_mult1_un54_sum_ac0_3_0_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001010110000"
        )
    port map (
            in0 => \N__14273\,
            in1 => \N__14350\,
            in2 => \N__13094\,
            in3 => \N__13090\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un4_haddress_if_m1_1_LC_6_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14351\,
            in1 => \_gnd_net_\,
            in2 => \N__13073\,
            in3 => \N__13821\,
            lcout => \this_vga_signals.if_m1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_1_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__14501\,
            in1 => \N__31014\,
            in2 => \N__13060\,
            in3 => \N__16169\,
            lcout => \this_vga_ramdac.N_3139_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_hcounter_d_cry_1_c_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15584\,
            in2 => \N__15538\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_2_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29783\,
            in1 => \N__13911\,
            in2 => \_gnd_net_\,
            in3 => \N__13211\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_1\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_3_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29787\,
            in1 => \N__13972\,
            in2 => \_gnd_net_\,
            in3 => \N__13208\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_2\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_4_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29784\,
            in1 => \N__13826\,
            in2 => \_gnd_net_\,
            in3 => \N__13205\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_3\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_5_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29788\,
            in1 => \N__14360\,
            in2 => \_gnd_net_\,
            in3 => \N__13202\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_4\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_6_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29785\,
            in1 => \N__14283\,
            in2 => \_gnd_net_\,
            in3 => \N__13199\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_6\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_5\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_7_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29789\,
            in1 => \N__14077\,
            in2 => \_gnd_net_\,
            in3 => \N__13196\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_7\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_6\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_8_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29786\,
            in1 => \N__14149\,
            in2 => \_gnd_net_\,
            in3 => \N__13193\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_8\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_hcounter_d_cry_7\,
            carryout => \this_vga_signals.un1_M_hcounter_d_cry_8\,
            clk => \N__39381\,
            ce => 'H',
            sr => \N__16289\
        );

    \this_vga_signals.M_hcounter_q_esr_9_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14216\,
            in2 => \_gnd_net_\,
            in3 => \N__13190\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39386\,
            ce => \N__16259\,
            sr => \N__16285\
        );

    \this_vga_signals.M_pcounter_q_0_e_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16313\,
            in1 => \N__16247\,
            in2 => \_gnd_net_\,
            in3 => \N__28615\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39393\,
            ce => \N__29792\,
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_13_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13334\,
            in2 => \_gnd_net_\,
            in3 => \N__23988\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_14_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23989\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13310\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_2_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23992\,
            in2 => \_gnd_net_\,
            in3 => \N__13541\,
            lcout => \this_ppu.oam_cache.N_823_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_5_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13583\,
            lcout => \this_ppu.oam_cache.N_820_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_7_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13277\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23993\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_8_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__23991\,
            in1 => \N__13253\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_9_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13232\,
            in2 => \_gnd_net_\,
            in3 => \N__23994\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_0_c_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23987\,
            in2 => \N__13449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_20_0_\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_LUT4_0_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13359\,
            in2 => \_gnd_net_\,
            in3 => \N__13214\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_0\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_LUT4_0_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13408\,
            in3 => \N__13484\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_1\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_LUT4_0_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13700\,
            in2 => \_gnd_net_\,
            in3 => \N__13481\,
            lcout => \this_ppu.un1_M_oam_cache_cnt_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_oam_cache_cnt_q_cry_2\,
            carryout => \this_ppu.un1_M_oam_cache_cnt_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__13475\,
            in1 => \N__21623\,
            in2 => \N__21524\,
            in3 => \N__13478\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39399\,
            ce => 'H',
            sr => \N__38962\
        );

    \this_ppu.M_state_q_ns_11_0__m71_i_o2_1_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13358\,
            in1 => \N__18247\,
            in2 => \N__13704\,
            in3 => \N__18407\,
            lcout => \this_ppu.m71_i_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m71_i_o2_0_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13442\,
            in1 => \N__18339\,
            in2 => \N__13407\,
            in3 => \N__18544\,
            lcout => OPEN,
            ltout => \this_ppu.m71_i_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m71_i_o2_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__18670\,
            in1 => \N__13474\,
            in2 => \N__13463\,
            in3 => \N__13460\,
            lcout => \this_ppu.N_796_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_cache_cnt_q_0_LC_7_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001001011010"
        )
    port map (
            in0 => \N__23983\,
            in1 => \N__21612\,
            in2 => \N__13450\,
            in3 => \N__21522\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39404\,
            ce => 'H',
            sr => \N__38959\
        );

    \this_ppu.M_oam_cache_cnt_q_2_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__13418\,
            in2 => \N__21622\,
            in3 => \N__13400\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39404\,
            ce => 'H',
            sr => \N__38959\
        );

    \this_ppu.M_oam_cache_cnt_q_1_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001001011010"
        )
    port map (
            in0 => \N__13360\,
            in1 => \N__21613\,
            in2 => \N__13376\,
            in3 => \N__21523\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39404\,
            ce => 'H',
            sr => \N__38959\
        );

    \this_ppu.M_oam_cache_cnt_q_3_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000111100"
        )
    port map (
            in0 => \N__21521\,
            in1 => \N__13715\,
            in2 => \N__13705\,
            in3 => \N__21620\,
            lcout => \this_ppu.M_oam_cache_cnt_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39404\,
            ce => 'H',
            sr => \N__38959\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_LC_7_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13604\,
            lcout => \this_ppu.oam_cache.N_826_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_1_LC_7_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23978\,
            in2 => \_gnd_net_\,
            in3 => \N__14018\,
            lcout => \this_ppu.oam_cache.N_824_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_4_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14036\,
            lcout => \this_ppu.oam_cache.N_821_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_3_LC_7_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23979\,
            in2 => \_gnd_net_\,
            in3 => \N__13502\,
            lcout => \this_ppu.oam_cache.N_822_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_6_LC_7_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13520\,
            lcout => \this_ppu.oam_cache.N_819_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_0_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23977\,
            in2 => \_gnd_net_\,
            in3 => \N__13562\,
            lcout => \this_ppu.oam_cache.N_825_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_state_q_7_i_a2_7_4_LC_7_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13597\,
            in1 => \N__13579\,
            in2 => \N__13561\,
            in3 => \N__13534\,
            lcout => \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_state_q_7_i_a2_7_3_LC_7_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13516\,
            in2 => \_gnd_net_\,
            in3 => \N__13498\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_state_q_7_i_a2_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_state_q_7_i_a2_7_LC_7_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__14032\,
            in1 => \N__14014\,
            in2 => \N__14000\,
            in3 => \N__13997\,
            lcout => \this_ppu.N_838_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m48_i_a2_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24050\,
            in2 => \_gnd_net_\,
            in3 => \N__21784\,
            lcout => \this_ppu.m48_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_11_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__21377\,
            in1 => \N__21722\,
            in2 => \_gnd_net_\,
            in3 => \N__36959\,
            lcout => \this_ppu.M_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_a2_3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18860\,
            lcout => OPEN,
            ltout => \this_ppu.m35_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_a2_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18240\,
            in1 => \N__18666\,
            in2 => \N__13991\,
            in3 => \N__16814\,
            lcout => \this_ppu.N_802\,
            ltout => \this_ppu.N_802_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_2_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__17090\,
            in1 => \_gnd_net_\,
            in2 => \N__13988\,
            in3 => \N__36960\,
            lcout => \this_ppu.M_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39357\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI3H6I_2_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13960\,
            in2 => \_gnd_net_\,
            in3 => \N__13900\,
            lcout => \this_vga_signals.un2_hsynclto3_1\,
            ltout => \this_vga_signals.un2_hsynclto3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_RNI58GD1_0_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__15559\,
            in1 => \N__15519\,
            in2 => \N__13853\,
            in3 => \N__13830\,
            lcout => \this_vga_signals.M_hcounter_d7lt7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_q_ret_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__30985\,
            in1 => \N__26491\,
            in2 => \N__13767\,
            in3 => \N__16159\,
            lcout => \this_vga_ramdac.M_this_vga_ramdac_en_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m10_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100101111"
        )
    port map (
            in0 => \N__14530\,
            in1 => \N__14609\,
            in2 => \N__14585\,
            in3 => \N__14560\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_2_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__30987\,
            in1 => \N__14422\,
            in2 => \N__14429\,
            in3 => \N__16158\,
            lcout => \this_vga_ramdac.N_3140_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m2_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__14559\,
            in2 => \_gnd_net_\,
            in3 => \N__14608\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.N_24_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_0_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__30986\,
            in1 => \N__14398\,
            in2 => \N__14408\,
            in3 => \N__16157\,
            lcout => \this_vga_ramdac.N_3138_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_6_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14387\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39366\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIVCD62_9_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__14370\,
            in1 => \N__14219\,
            in2 => \N__14306\,
            in3 => \N__14294\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_864_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNITLAV2_9_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__14220\,
            in1 => \N__14165\,
            in2 => \N__14108\,
            in3 => \N__14093\,
            lcout => \this_vga_signals.M_hcounter_d7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m16_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110010111"
        )
    port map (
            in0 => \N__14580\,
            in1 => \N__14557\,
            in2 => \N__14533\,
            in3 => \N__14606\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_3_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__14644\,
            in1 => \N__30988\,
            in2 => \N__14657\,
            in3 => \N__16164\,
            lcout => \this_vga_ramdac.N_3141_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m19_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100100101011"
        )
    port map (
            in0 => \N__14581\,
            in1 => \N__14558\,
            in2 => \N__14534\,
            in3 => \N__14607\,
            lcout => OPEN,
            ltout => \this_vga_ramdac.m19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_4_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__14620\,
            in1 => \N__30989\,
            in2 => \N__14633\,
            in3 => \N__16165\,
            lcout => \this_vga_ramdac.N_3142_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39374\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m22_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100011001"
        )
    port map (
            in0 => \N__14579\,
            in1 => \N__14556\,
            in2 => \N__14532\,
            in3 => \N__14605\,
            lcout => \this_vga_ramdac.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_5_0__m6_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000111111"
        )
    port map (
            in0 => \N__14604\,
            in1 => \N__14578\,
            in2 => \N__14561\,
            in3 => \N__14520\,
            lcout => \this_vga_ramdac.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNID8M7_17_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14477\,
            lcout => \this_ppu.M_oam_cache_read_data_i_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_17_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14489\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_16_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14471\,
            lcout => \this_ppu.M_oam_cache_read_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_ramdac.M_this_rgb_d_3_0_dreg_5_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__14459\,
            in1 => \N__30991\,
            in2 => \N__14446\,
            in3 => \N__16160\,
            lcout => \this_vga_ramdac.N_3143_reto\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_1_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001100010"
        )
    port map (
            in0 => \N__16243\,
            in1 => \N__29774\,
            in2 => \N__16219\,
            in3 => \N__28586\,
            lcout => \this_vga_signals.M_pcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_18_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIC31GS_2_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__18408\,
            in1 => \N__18800\,
            in2 => \N__18350\,
            in3 => \N__18452\,
            lcout => \this_ppu.N_777_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIKRNBS_1_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18409\,
            in1 => \N__18798\,
            in2 => \_gnd_net_\,
            in3 => \N__18451\,
            lcout => \this_ppu.N_776_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14774\,
            in1 => \N__14762\,
            in2 => \N__14786\,
            in3 => \N__14804\,
            lcout => \this_ppu.N_932_0\,
            ltout => \this_ppu.N_932_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_0_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110001"
        )
    port map (
            in0 => \N__17258\,
            in1 => \N__23849\,
            in2 => \N__14705\,
            in3 => \N__14677\,
            lcout => \this_ppu.un1_M_state_q_7_i_0_0\,
            ltout => \this_ppu.un1_M_state_q_7_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNITKE7S_0_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000100010"
        )
    port map (
            in0 => \N__18799\,
            in1 => \N__18540\,
            in2 => \N__14702\,
            in3 => \N__18578\,
            lcout => \this_ppu.N_775_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_3_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__17259\,
            in1 => \N__14684\,
            in2 => \_gnd_net_\,
            in3 => \N__14678\,
            lcout => \this_ppu.M_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39389\,
            ce => 'H',
            sr => \N__36831\
        );

    \this_ppu.un1_oam_data_1_cry_0_c_inv_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14663\,
            in2 => \N__22742\,
            in3 => \N__23482\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_9_21_0_\,
            carryout => \this_ppu.un1_oam_data_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_1_c_inv_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14816\,
            in2 => \N__22694\,
            in3 => \N__23437\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_17\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_0\,
            carryout => \this_ppu.un1_oam_data_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_2_c_inv_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14810\,
            in2 => \N__22652\,
            in3 => \N__23398\,
            lcout => \this_ppu.M_this_oam_ram_read_data_i_18\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_1\,
            carryout => \this_ppu.un1_oam_data_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m28_e_i_o2_0_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000001"
        )
    port map (
            in0 => \N__14795\,
            in1 => \N__15116\,
            in2 => \N__22606\,
            in3 => \N__14798\,
            lcout => \this_ppu.m28_e_i_o2_0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_2\,
            carryout => \this_ppu.un1_oam_data_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_3_c_RNIT7ID_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15482\,
            in2 => \N__22555\,
            in3 => \N__14789\,
            lcout => \this_ppu.un1_oam_data_1_cry_3_c_RNIT7IDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_3\,
            carryout => \this_ppu.un1_oam_data_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJD_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14996\,
            in2 => \N__22495\,
            in3 => \N__14777\,
            lcout => \this_ppu.un1_oam_data_1_cry_4_c_RNIVAJDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_4\,
            carryout => \this_ppu.un1_oam_data_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKD_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14954\,
            in2 => \N__22438\,
            in3 => \N__14768\,
            lcout => \this_ppu.un1_oam_data_1_cry_5_c_RNI1EKDZ0\,
            ltout => OPEN,
            carryin => \this_ppu.un1_oam_data_1_cry_5\,
            carryout => \this_ppu.un1_oam_data_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLD_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__23296\,
            in2 => \_gnd_net_\,
            in3 => \N__14765\,
            lcout => \this_ppu.un1_oam_data_1_cry_6_c_RNI3HLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_4_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15017\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_5_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23885\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_2_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14971\,
            lcout => \M_this_oam_ram_read_data_i_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_6_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23886\,
            in2 => \_gnd_net_\,
            in3 => \N__14948\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_7_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23883\,
            in2 => \_gnd_net_\,
            in3 => \N__14918\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_8_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14891\,
            in2 => \_gnd_net_\,
            in3 => \N__23887\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_9_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23882\,
            in2 => \_gnd_net_\,
            in3 => \N__14870\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_6_LC_9_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37389\,
            lcout => \M_this_data_tmp_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39420\,
            ce => \N__23620\,
            sr => \N__36841\
        );

    \M_this_data_tmp_q_esr_3_LC_9_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39420\,
            ce => \N__23620\,
            sr => \N__36841\
        );

    \this_start_data_delay.M_last_q_RNIPR151_LC_9_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19370\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16661\,
            lcout => \M_this_oam_ram_write_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_13_LC_9_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14840\,
            in2 => \_gnd_net_\,
            in3 => \N__23972\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOQ151_LC_9_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17153\,
            in2 => \_gnd_net_\,
            in3 => \N__19373\,
            lcout => \M_this_oam_ram_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIQS151_LC_9_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17162\,
            lcout => \M_this_oam_ram_write_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNITV151_LC_9_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21881\,
            in2 => \_gnd_net_\,
            in3 => \N__19369\,
            lcout => \M_this_oam_ram_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_14_LC_9_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23971\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15062\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICRDD1_LC_9_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16667\,
            in2 => \_gnd_net_\,
            in3 => \N__19372\,
            lcout => \M_this_oam_ram_write_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI7MDD1_LC_9_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15032\,
            lcout => \M_this_oam_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_1_LC_9_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15013\,
            lcout => \M_this_oam_ram_read_data_i_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIAPDD1_LC_9_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14987\,
            lcout => \M_this_oam_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI9ODD1_LC_9_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19376\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16619\,
            lcout => \M_this_oam_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBQDD1_LC_9_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16625\,
            in2 => \_gnd_net_\,
            in3 => \N__19374\,
            lcout => \M_this_oam_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_11_LC_9_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15197\,
            in2 => \_gnd_net_\,
            in3 => \N__23973\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_12_LC_9_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15176\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIRT151_LC_9_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19365\,
            in2 => \_gnd_net_\,
            in3 => \N__16607\,
            lcout => \M_this_oam_ram_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOR251_LC_9_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19378\,
            lcout => \M_this_oam_ram_write_data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_2_LC_9_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23976\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_LC_9_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15127\,
            lcout => \M_this_oam_ram_read_data_i_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_3_LC_9_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23974\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_oam_ram.mem_mem_0_1_RNITG75_0_LC_9_30_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15493\,
            lcout => \M_this_oam_ram_read_data_i_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI43IG1_LC_9_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19380\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37853\,
            lcout => \M_this_oam_ram_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI76IG1_LC_9_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37397\,
            in2 => \_gnd_net_\,
            in3 => \N__19382\,
            lcout => \M_this_oam_ram_write_data_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNISU151_LC_9_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19383\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17540\,
            lcout => \M_this_oam_ram_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI65IG1_LC_9_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19381\,
            lcout => \M_this_oam_ram_write_data_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI10IG1_LC_9_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => \M_this_oam_ram_write_data_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dma_0_sbtinv_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => dma_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_7_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15239\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_3_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15224\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_4_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15635\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39323\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__15620\,
            in1 => \N__15610\,
            in2 => \_gnd_net_\,
            in3 => \N__36928\,
            lcout => \this_pixel_clk_M_counter_q_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.G_424_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15619\,
            in1 => \N__15609\,
            in2 => \_gnd_net_\,
            in3 => \N__36927\,
            lcout => \this_vga_signals.GZ0Z_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_pixel_clk.M_counter_q_0_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15611\,
            lcout => \this_pixel_clk_M_counter_q_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39339\,
            ce => 'H',
            sr => \N__36825\
        );

    \this_vga_signals.M_hcounter_q_1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15529\,
            in2 => \N__29779\,
            in3 => \N__15577\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39350\,
            ce => 'H',
            sr => \N__16278\
        );

    \this_vga_signals.M_hcounter_q_0_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__15530\,
            in1 => \N__29743\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_hcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39350\,
            ce => 'H',
            sr => \N__16278\
        );

    \this_ppu.oam_cache.read_data_RNI61M7_10_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16364\,
            lcout => \this_ppu.M_oam_cache_read_data_i_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_e_RNICJLB4_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16215\,
            in1 => \N__29731\,
            in2 => \_gnd_net_\,
            in3 => \N__16295\,
            lcout => \N_3_0\,
            ltout => \N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_2_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15497\,
            in3 => \N__16193\,
            lcout => \M_this_vga_signals_pixel_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_pcounter_q_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39358\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_ret_RNITMRI3_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16306\,
            in1 => \N__16241\,
            in2 => \_gnd_net_\,
            in3 => \N__28567\,
            lcout => \this_vga_signals.M_pcounter_q_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNIIG783_9_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29732\,
            lcout => \this_vga_signals.N_1188_1\,
            ltout => \this_vga_signals.N_1188_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_hcounter_q_esr_RNO_0_9_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29734\,
            in1 => \_gnd_net_\,
            in2 => \N__16262\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.N_933_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_pcounter_q_0_RNI38654_1_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011001100"
        )
    port map (
            in0 => \N__28568\,
            in1 => \N__16242\,
            in2 => \N__16220\,
            in3 => \N__29733\,
            lcout => \N_2_0\,
            ltout => \N_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__G_462_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16187\,
            in2 => \N__16181\,
            in3 => \N__16177\,
            lcout => \G_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_y_cry_0_c_inv_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17512\,
            in1 => \N__22741\,
            in2 => \N__16127\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_oam_cache_read_data_i_16\,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \this_ppu.offset_y_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_y_cry_0_c_RNIVBJT1_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100110011100"
        )
    port map (
            in0 => \N__32689\,
            in1 => \N__22693\,
            in2 => \N__16118\,
            in3 => \N__15905\,
            lcout => \M_this_ppu_spr_addr_4\,
            ltout => OPEN,
            carryin => \this_ppu.offset_y_cry_0\,
            carryout => \this_ppu.offset_y_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI2GKT1_18_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011001001"
        )
    port map (
            in0 => \N__15902\,
            in1 => \N__22651\,
            in2 => \N__32705\,
            in3 => \N__15896\,
            lcout => \M_this_ppu_spr_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_10_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16373\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m18_i_m2_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__17263\,
            in1 => \N__21568\,
            in2 => \N__18841\,
            in3 => \N__21505\,
            lcout => OPEN,
            ltout => \this_ppu.N_836_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_1_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__31012\,
            in1 => \_gnd_net_\,
            in2 => \N__16355\,
            in3 => \N__18468\,
            lcout => \this_ppu.M_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m13_0_a2_0_0_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__21785\,
            in1 => \N__21721\,
            in2 => \_gnd_net_\,
            in3 => \N__21567\,
            lcout => \this_ppu.m13_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_9_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_M_this_warmup_d_cry_1_c_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17071\,
            in2 => \N__17060\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \un1_M_this_warmup_d_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_warmup_q_2_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16340\,
            in2 => \_gnd_net_\,
            in3 => \N__16334\,
            lcout => \M_this_warmup_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_1\,
            carryout => \un1_M_this_warmup_d_cry_2\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_3_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16331\,
            in2 => \_gnd_net_\,
            in3 => \N__16325\,
            lcout => \M_this_warmup_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_2\,
            carryout => \un1_M_this_warmup_d_cry_3\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_4_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16322\,
            in2 => \_gnd_net_\,
            in3 => \N__16316\,
            lcout => \M_this_warmup_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_3\,
            carryout => \un1_M_this_warmup_d_cry_4\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_5_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16451\,
            in2 => \_gnd_net_\,
            in3 => \N__16445\,
            lcout => \M_this_warmup_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_4\,
            carryout => \un1_M_this_warmup_d_cry_5\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_6_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16442\,
            in2 => \_gnd_net_\,
            in3 => \N__16436\,
            lcout => \M_this_warmup_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_5\,
            carryout => \un1_M_this_warmup_d_cry_6\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_7_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16433\,
            in2 => \_gnd_net_\,
            in3 => \N__16427\,
            lcout => \M_this_warmup_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_6\,
            carryout => \un1_M_this_warmup_d_cry_7\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_8_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16424\,
            in2 => \_gnd_net_\,
            in3 => \N__16418\,
            lcout => \M_this_warmup_qZ0Z_8\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_7\,
            carryout => \un1_M_this_warmup_d_cry_8\,
            clk => \N__39375\,
            ce => 'H',
            sr => \N__36829\
        );

    \M_this_warmup_q_9_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16415\,
            in2 => \_gnd_net_\,
            in3 => \N__16409\,
            lcout => \M_this_warmup_qZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \un1_M_this_warmup_d_cry_9\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_10_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16406\,
            in2 => \_gnd_net_\,
            in3 => \N__16400\,
            lcout => \M_this_warmup_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_9\,
            carryout => \un1_M_this_warmup_d_cry_10\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_11_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \_gnd_net_\,
            in3 => \N__16391\,
            lcout => \M_this_warmup_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_10\,
            carryout => \un1_M_this_warmup_d_cry_11\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_12_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16388\,
            in2 => \_gnd_net_\,
            in3 => \N__16382\,
            lcout => \M_this_warmup_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_11\,
            carryout => \un1_M_this_warmup_d_cry_12\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_13_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16379\,
            in2 => \_gnd_net_\,
            in3 => \N__16526\,
            lcout => \M_this_warmup_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_12\,
            carryout => \un1_M_this_warmup_d_cry_13\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_14_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16523\,
            in2 => \_gnd_net_\,
            in3 => \N__16517\,
            lcout => \M_this_warmup_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_13\,
            carryout => \un1_M_this_warmup_d_cry_14\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_15_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16514\,
            in2 => \_gnd_net_\,
            in3 => \N__16508\,
            lcout => \M_this_warmup_qZ0Z_15\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_14\,
            carryout => \un1_M_this_warmup_d_cry_15\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_16_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16505\,
            in2 => \_gnd_net_\,
            in3 => \N__16499\,
            lcout => \M_this_warmup_qZ0Z_16\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_15\,
            carryout => \un1_M_this_warmup_d_cry_16\,
            clk => \N__39383\,
            ce => 'H',
            sr => \N__36830\
        );

    \M_this_warmup_q_17_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16496\,
            in2 => \_gnd_net_\,
            in3 => \N__16490\,
            lcout => \M_this_warmup_qZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \un1_M_this_warmup_d_cry_17\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_18_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16487\,
            in2 => \_gnd_net_\,
            in3 => \N__16481\,
            lcout => \M_this_warmup_qZ0Z_18\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_17\,
            carryout => \un1_M_this_warmup_d_cry_18\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_19_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16478\,
            in2 => \_gnd_net_\,
            in3 => \N__16472\,
            lcout => \M_this_warmup_qZ0Z_19\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_18\,
            carryout => \un1_M_this_warmup_d_cry_19\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_20_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16469\,
            in2 => \_gnd_net_\,
            in3 => \N__16463\,
            lcout => \M_this_warmup_qZ0Z_20\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_19\,
            carryout => \un1_M_this_warmup_d_cry_20\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_21_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16460\,
            in2 => \_gnd_net_\,
            in3 => \N__16454\,
            lcout => \M_this_warmup_qZ0Z_21\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_20\,
            carryout => \un1_M_this_warmup_d_cry_21\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_22_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16592\,
            in2 => \_gnd_net_\,
            in3 => \N__16586\,
            lcout => \M_this_warmup_qZ0Z_22\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_21\,
            carryout => \un1_M_this_warmup_d_cry_22\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_23_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16583\,
            in2 => \_gnd_net_\,
            in3 => \N__16577\,
            lcout => \M_this_warmup_qZ0Z_23\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_22\,
            carryout => \un1_M_this_warmup_d_cry_23\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_24_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16574\,
            in2 => \_gnd_net_\,
            in3 => \N__16568\,
            lcout => \M_this_warmup_qZ0Z_24\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_23\,
            carryout => \un1_M_this_warmup_d_cry_24\,
            clk => \N__39390\,
            ce => 'H',
            sr => \N__36832\
        );

    \M_this_warmup_q_25_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16565\,
            in2 => \_gnd_net_\,
            in3 => \N__16559\,
            lcout => \M_this_warmup_qZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \un1_M_this_warmup_d_cry_25\,
            clk => \N__39394\,
            ce => 'H',
            sr => \N__36833\
        );

    \M_this_warmup_q_26_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16556\,
            in2 => \_gnd_net_\,
            in3 => \N__16550\,
            lcout => \M_this_warmup_qZ0Z_26\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_25\,
            carryout => \un1_M_this_warmup_d_cry_26\,
            clk => \N__39394\,
            ce => 'H',
            sr => \N__36833\
        );

    \M_this_warmup_q_27_LC_10_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16547\,
            in2 => \_gnd_net_\,
            in3 => \N__16541\,
            lcout => \M_this_warmup_qZ0Z_27\,
            ltout => OPEN,
            carryin => \un1_M_this_warmup_d_cry_26\,
            carryout => \un1_M_this_warmup_d_cry_27\,
            clk => \N__39394\,
            ce => 'H',
            sr => \N__36833\
        );

    \M_this_warmup_q_28_LC_10_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16534\,
            in2 => \_gnd_net_\,
            in3 => \N__16538\,
            lcout => \M_this_warmup_qZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39394\,
            ce => 'H',
            sr => \N__36833\
        );

    \M_this_status_flags_q_0_LC_10_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18831\,
            lcout => \M_this_status_flags_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39394\,
            ce => 'H',
            sr => \N__36833\
        );

    \M_this_data_tmp_q_esr_8_LC_10_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38103\,
            lcout => \M_this_data_tmp_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39411\,
            ce => \N__19426\,
            sr => \N__36837\
        );

    \M_this_data_tmp_q_esr_14_LC_10_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37388\,
            lcout => \M_this_data_tmp_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39411\,
            ce => \N__19426\,
            sr => \N__36837\
        );

    \M_this_data_tmp_q_esr_10_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39411\,
            ce => \N__19426\,
            sr => \N__36837\
        );

    \this_start_data_delay.M_last_q_RNILN151_LC_10_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16655\,
            in2 => \_gnd_net_\,
            in3 => \N__19328\,
            lcout => \M_this_oam_ram_write_data_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINP151_LC_10_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17168\,
            in2 => \_gnd_net_\,
            in3 => \N__19327\,
            lcout => \M_this_oam_ram_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_7_LC_10_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38729\,
            lcout => \M_this_data_tmp_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39421\,
            ce => \N__23621\,
            sr => \N__36842\
        );

    \M_this_data_tmp_q_esr_5_LC_10_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39421\,
            ce => \N__23621\,
            sr => \N__36842\
        );

    \M_this_data_tmp_q_esr_22_LC_10_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39427\,
            ce => \N__21851\,
            sr => \N__36845\
        );

    \M_this_data_tmp_q_esr_16_LC_10_30_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38101\,
            lcout => \M_this_data_tmp_qZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39427\,
            ce => \N__21851\,
            sr => \N__36845\
        );

    \this_start_data_delay.M_last_q_RNI87IG1_LC_10_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19364\,
            lcout => \M_this_oam_ram_write_data_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINQ251_LC_10_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19363\,
            in1 => \N__19844\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_write_data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIPS251_LC_10_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19362\,
            in2 => \_gnd_net_\,
            in3 => \N__17774\,
            lcout => \M_this_oam_ram_write_data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_wclke_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__32222\,
            in1 => \N__32126\,
            in2 => \N__32036\,
            in3 => \N__31919\,
            lcout => \this_spr_ram.mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_wclke_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__32218\,
            in1 => \N__32125\,
            in2 => \N__32032\,
            in3 => \N__31914\,
            lcout => \this_spr_ram.mem_WE_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_5_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16736\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39310\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_7_0_wclke_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32213\,
            in1 => \N__32118\,
            in2 => \N__32030\,
            in3 => \N__31898\,
            lcout => \this_spr_ram.mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_34_i_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__17892\,
            in1 => \N__22136\,
            in2 => \N__18752\,
            in3 => \N__19628\,
            lcout => \N_34_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_14_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16682\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI3UQE7_4_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__21780\,
            in1 => \N__21579\,
            in2 => \N__21374\,
            in3 => \N__21519\,
            lcout => \this_ppu.M_oam_curr_qc_0_1\,
            ltout => \this_ppu.M_oam_curr_qc_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_3_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18223\,
            in2 => \N__16817\,
            in3 => \N__18274\,
            lcout => \M_this_ppu_oam_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39324\,
            ce => 'H',
            sr => \N__38963\
        );

    \this_ppu.M_oam_curr_q_4_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110000000000"
        )
    port map (
            in0 => \N__18275\,
            in1 => \N__18650\,
            in2 => \N__18236\,
            in3 => \N__18889\,
            lcout => \M_this_ppu_oam_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39324\,
            ce => 'H',
            sr => \N__38963\
        );

    \this_ppu.M_oam_curr_q_2_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100011000000"
        )
    port map (
            in0 => \N__18388\,
            in1 => \N__18888\,
            in2 => \N__18317\,
            in3 => \N__18445\,
            lcout => \M_this_ppu_oam_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39324\,
            ce => 'H',
            sr => \N__38963\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_a2_4_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18387\,
            in1 => \N__18304\,
            in2 => \N__18926\,
            in3 => \N__18517\,
            lcout => \this_ppu.m35_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_1_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18392\,
            in1 => \N__18885\,
            in2 => \_gnd_net_\,
            in3 => \N__18444\,
            lcout => \M_this_ppu_oam_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39332\,
            ce => 'H',
            sr => \N__38960\
        );

    \this_ppu.M_oam_curr_q_0_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001000001010"
        )
    port map (
            in0 => \N__18886\,
            in1 => \N__18570\,
            in2 => \N__18533\,
            in3 => \N__18476\,
            lcout => \M_this_ppu_oam_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39332\,
            ce => 'H',
            sr => \N__38960\
        );

    \this_ppu.M_screen_x_q_1_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__17143\,
            in1 => \N__16965\,
            in2 => \N__16942\,
            in3 => \N__16862\,
            lcout => \M_this_ppu_vram_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_5_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__17016\,
            in1 => \N__17141\,
            in2 => \_gnd_net_\,
            in3 => \N__17036\,
            lcout => \M_this_ppu_vram_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_0_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__22269\,
            in1 => \N__30900\,
            in2 => \N__16941\,
            in3 => \N__16861\,
            lcout => \M_this_ppu_vram_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIB9B9C_11_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111110"
        )
    port map (
            in0 => \N__20971\,
            in1 => \N__21114\,
            in2 => \N__21166\,
            in3 => \N__21188\,
            lcout => \this_ppu.N_827_0\,
            ltout => \this_ppu.N_827_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNIM77RC_1_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16964\,
            in2 => \N__17042\,
            in3 => \N__16927\,
            lcout => \this_ppu.un1_M_screen_x_q_c2\,
            ltout => \this_ppu.un1_M_screen_x_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNIUC1MD_4_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16833\,
            in1 => \N__16883\,
            in2 => \N__17039\,
            in3 => \N__17880\,
            lcout => \this_ppu.un1_M_screen_x_q_c5\,
            ltout => \this_ppu.un1_M_screen_x_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010001000"
        )
    port map (
            in0 => \N__17142\,
            in1 => \N__16993\,
            in2 => \N__17030\,
            in3 => \N__17017\,
            lcout => \M_this_ppu_vram_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_2_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__30899\,
            in1 => \N__22270\,
            in2 => \N__16896\,
            in3 => \N__16982\,
            lcout => \M_this_ppu_vram_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_RNID854D_1_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16966\,
            in1 => \N__16928\,
            in2 => \N__16900\,
            in3 => \N__16860\,
            lcout => \this_ppu.un1_M_screen_x_q_c3\,
            ltout => \this_ppu.un1_M_screen_x_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_4_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110000000000"
        )
    port map (
            in0 => \N__17885\,
            in1 => \N__16834\,
            in2 => \N__16847\,
            in3 => \N__17144\,
            lcout => \M_this_ppu_vram_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_6_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19160\,
            in1 => \N__21440\,
            in2 => \N__30932\,
            in3 => \N__19025\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_0_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__19001\,
            in1 => \N__28654\,
            in2 => \_gnd_net_\,
            in3 => \N__28596\,
            lcout => \this_vga_signals.i22_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIGL6V4_0_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__30894\,
            in1 => \N__21569\,
            in2 => \_gnd_net_\,
            in3 => \N__21506\,
            lcout => \this_ppu.N_1210_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_x_q_3_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__17884\,
            in1 => \N__30895\,
            in2 => \N__22274\,
            in3 => \N__17126\,
            lcout => \M_this_ppu_vram_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39351\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21439\,
            in1 => \N__21209\,
            in2 => \N__31019\,
            in3 => \N__19159\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_13_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17120\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_12_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17111\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m13_0_a2_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21647\,
            in1 => \N__21570\,
            in2 => \_gnd_net_\,
            in3 => \N__21504\,
            lcout => OPEN,
            ltout => \this_ppu.N_844_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_0_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21373\,
            in1 => \N__17102\,
            in2 => \N__17093\,
            in3 => \N__31011\,
            lcout => \this_ppu.M_state_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39359\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIRJK11_1_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21113\,
            in1 => \N__23951\,
            in2 => \N__20977\,
            in3 => \N__17083\,
            lcout => \this_ppu.un1_M_pixel_cnt_d_1_sqmuxa_0_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_warmup_q_1_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__17059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17072\,
            lcout => \M_this_warmup_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39368\,
            ce => 'H',
            sr => \N__36828\
        );

    \M_this_warmup_q_0_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17058\,
            lcout => \M_this_warmup_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39368\,
            ce => 'H',
            sr => \N__36828\
        );

    \this_ppu.oam_cache.read_data_RNIUU07_9_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17528\,
            lcout => \this_ppu.M_oam_cache_read_data_i_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI62LG1_16_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__32670\,
            in1 => \N__17522\,
            in2 => \_gnd_net_\,
            in3 => \N__22737\,
            lcout => \M_this_ppu_spr_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI41OT_2_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21714\,
            in1 => \N__20978\,
            in2 => \N__17270\,
            in3 => \N__23955\,
            lcout => \this_ppu_N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_6_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17214\,
            in1 => \N__25212\,
            in2 => \_gnd_net_\,
            in3 => \N__19435\,
            lcout => \M_this_oam_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39405\,
            ce => 'H',
            sr => \N__38952\
        );

    \M_this_oam_address_q_7_LC_11_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__19436\,
            in1 => \N__17182\,
            in2 => \N__25217\,
            in3 => \N__17215\,
            lcout => \M_this_oam_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39405\,
            ce => 'H',
            sr => \N__38952\
        );

    \M_this_data_tmp_q_esr_20_LC_11_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37466\,
            lcout => \M_this_data_tmp_qZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39408\,
            ce => \N__21824\,
            sr => \N__36835\
        );

    \M_this_data_tmp_q_esr_12_LC_11_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37506\,
            lcout => \M_this_data_tmp_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39412\,
            ce => \N__19427\,
            sr => \N__36838\
        );

    \M_this_data_tmp_q_esr_15_LC_11_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38768\,
            lcout => \M_this_data_tmp_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39412\,
            ce => \N__19427\,
            sr => \N__36838\
        );

    \M_this_data_tmp_q_esr_13_LC_11_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38917\,
            lcout => \M_this_data_tmp_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39412\,
            ce => \N__19427\,
            sr => \N__36838\
        );

    \M_this_data_tmp_q_esr_11_LC_11_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39412\,
            ce => \N__19427\,
            sr => \N__36838\
        );

    \M_this_data_tmp_q_esr_9_LC_11_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37735\,
            lcout => \M_this_data_tmp_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39412\,
            ce => \N__19427\,
            sr => \N__36838\
        );

    \this_start_data_delay.M_last_q_RNI5KDD1_LC_11_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21869\,
            lcout => \M_this_oam_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIMP251_LC_11_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19297\,
            in2 => \_gnd_net_\,
            in3 => \N__17615\,
            lcout => \M_this_oam_ram_write_data_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI6LDD1_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19850\,
            lcout => \M_this_oam_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIDSDD1_LC_11_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19301\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17582\,
            lcout => \M_this_oam_ram_write_data_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI8NDD1_LC_11_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19296\,
            in2 => \_gnd_net_\,
            in3 => \N__19208\,
            lcout => \M_this_oam_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIMO151_LC_11_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19300\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17555\,
            lcout => \M_this_oam_ram_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_17_LC_11_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37734\,
            lcout => \M_this_data_tmp_qZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39422\,
            ce => \N__21850\,
            sr => \N__36843\
        );

    \M_this_data_tmp_q_esr_23_LC_11_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38769\,
            lcout => \M_this_data_tmp_qZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39422\,
            ce => \N__21850\,
            sr => \N__36843\
        );

    \this_start_data_delay.M_last_q_RNIU0251_LC_11_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21860\,
            in2 => \_gnd_net_\,
            in3 => \N__19384\,
            lcout => \M_this_oam_ram_write_data_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI54IG1_LC_11_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19386\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37507\,
            lcout => \M_this_oam_ram_write_data_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI21IG1_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37715\,
            in2 => \_gnd_net_\,
            in3 => \N__19385\,
            lcout => \M_this_oam_ram_write_data_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_0_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20825\,
            in1 => \N__17738\,
            in2 => \_gnd_net_\,
            in3 => \N__17723\,
            lcout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_0_12_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__19925\,
            in1 => \N__17936\,
            in2 => \N__19693\,
            in3 => \N__17711\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_0_11_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__19926\,
            in1 => \N__17633\,
            in2 => \N__17705\,
            in3 => \N__17672\,
            lcout => \M_this_spr_ram_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17702\,
            in1 => \N__17684\,
            in2 => \_gnd_net_\,
            in3 => \N__20839\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20840\,
            in1 => \N__17666\,
            in2 => \_gnd_net_\,
            in3 => \N__17651\,
            lcout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_0_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20826\,
            in1 => \N__17972\,
            in2 => \_gnd_net_\,
            in3 => \N__17954\,
            lcout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20827\,
            in1 => \N__17930\,
            in2 => \_gnd_net_\,
            in3 => \N__17915\,
            lcout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_12_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000011111"
        )
    port map (
            in0 => \N__19906\,
            in1 => \N__19967\,
            in2 => \N__19694\,
            in3 => \N__17903\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.m21_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17896\,
            in2 => \_gnd_net_\,
            in3 => \N__22135\,
            lcout => \this_vga_signals.N_22_0\,
            ltout => \this_vga_signals.N_22_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_856_i_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000100"
        )
    port map (
            in0 => \N__18748\,
            in1 => \N__22075\,
            in2 => \N__17849\,
            in3 => \N__18611\,
            lcout => \N_856_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17831\,
            in1 => \N__17813\,
            in2 => \_gnd_net_\,
            in3 => \N__20863\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_11_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__20780\,
            in1 => \N__19910\,
            in2 => \N__17798\,
            in3 => \N__17795\,
            lcout => \M_this_spr_ram_read_data_3\,
            ltout => \M_this_spr_ram_read_data_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_25_0_i_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__18747\,
            in1 => \N__18706\,
            in2 => \N__17789\,
            in3 => \N__22361\,
            lcout => \N_25_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIA5M7_14_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18161\,
            lcout => \this_ppu.M_oam_cache_read_data_i_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_1_RNIM6VF_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20852\,
            in1 => \N__18155\,
            in2 => \_gnd_net_\,
            in3 => \N__18137\,
            lcout => \this_spr_ram.mem_mem_0_1_RNIM6VFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNII6H51_6_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21163\,
            in1 => \N__20767\,
            in2 => \N__21778\,
            in3 => \N__22042\,
            lcout => \this_ppu.M_state_q_inv_1\,
            ltout => \this_ppu.M_state_q_inv_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_12_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18125\,
            in2 => \N__18113\,
            in3 => \N__18110\,
            lcout => \this_spr_ram.mem_radregZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39311\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_5_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__18571\,
            in1 => \N__21376\,
            in2 => \N__18089\,
            in3 => \N__30983\,
            lcout => \this_ppu.M_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39317\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_1_RNIOA1G_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18077\,
            in1 => \N__18059\,
            in2 => \_gnd_net_\,
            in3 => \N__20865\,
            lcout => \this_spr_ram.mem_mem_1_1_RNIOA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20866\,
            in1 => \N__18044\,
            in2 => \_gnd_net_\,
            in3 => \N__18029\,
            lcout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18011\,
            in1 => \N__20864\,
            in2 => \_gnd_net_\,
            in3 => \N__17993\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNITCNI1_0_12_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__19915\,
            in1 => \N__19682\,
            in2 => \N__17981\,
            in3 => \N__17978\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNINL8S2_0_11_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__19927\,
            in1 => \N__18767\,
            in2 => \N__18761\,
            in3 => \N__18758\,
            lcout => \M_this_spr_ram_read_data_2\,
            ltout => \M_this_spr_ram_read_data_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.N_28_0_i_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__18746\,
            in1 => \N__18710\,
            in2 => \N__18695\,
            in3 => \N__22397\,
            lcout => \N_28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIGIC2L_4_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18646\,
            in1 => \N__18221\,
            in2 => \_gnd_net_\,
            in3 => \N__18273\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_d25_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18617\,
            in1 => \N__18610\,
            in2 => \N__18596\,
            in3 => \N__19627\,
            lcout => \this_ppu.M_oam_curr_dZ0Z25\,
            ltout => \this_ppu.M_oam_curr_dZ0Z25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIQ09CG_6_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__22041\,
            in1 => \N__21165\,
            in2 => \N__18581\,
            in3 => \N__22015\,
            lcout => \this_ppu.N_834_0\,
            ltout => \this_ppu.N_834_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNIEH7HK_0_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18513\,
            in2 => \N__18479\,
            in3 => \N__18475\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c1\,
            ltout => \this_ppu.un1_M_oam_curr_q_1_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNITVPPK_2_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__18386\,
            in1 => \_gnd_net_\,
            in2 => \N__18353\,
            in3 => \N__18303\,
            lcout => \this_ppu.un1_M_oam_curr_q_1_c3\,
            ltout => \this_ppu.un1_M_oam_curr_q_1_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_RNI5CAKS_3_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__18222\,
            in1 => \_gnd_net_\,
            in2 => \N__18188\,
            in3 => \N__18787\,
            lcout => \this_ppu.N_778_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_oam_curr_q_5_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__18927\,
            in1 => \N__18887\,
            in2 => \_gnd_net_\,
            in3 => \N__18955\,
            lcout => \M_this_ppu_oam_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39325\,
            ce => 'H',
            sr => \N__38957\
        );

    \this_ppu.M_oam_curr_q_6_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110000000000"
        )
    port map (
            in0 => \N__18956\,
            in1 => \N__18859\,
            in2 => \N__18928\,
            in3 => \N__18890\,
            lcout => \this_ppu.M_oam_curr_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39325\,
            ce => 'H',
            sr => \N__38957\
        );

    \this_ppu.M_state_q_7_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30990\,
            in2 => \_gnd_net_\,
            in3 => \N__22019\,
            lcout => \this_ppu.M_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_10_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000010"
        )
    port map (
            in0 => \N__22250\,
            in1 => \N__18845\,
            in2 => \N__36963\,
            in3 => \N__20976\,
            lcout => \this_ppu.M_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_15_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18812\,
            lcout => \this_ppu.M_oam_cache_read_data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39333\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIF37M7_4_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__21779\,
            in1 => \N__36929\,
            in2 => \N__21359\,
            in3 => \N__22249\,
            lcout => \this_ppu.N_784_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNO_0_1_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18979\,
            in1 => \N__28655\,
            in2 => \_gnd_net_\,
            in3 => \N__28612\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_1_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010011001100"
        )
    port map (
            in0 => \N__28614\,
            in1 => \N__19000\,
            in2 => \N__18776\,
            in3 => \N__29778\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI94M7_13_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18773\,
            lcout => \this_ppu.M_oam_cache_read_data_i_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m9_0_a2_5_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19090\,
            in1 => \N__19066\,
            in2 => \N__19042\,
            in3 => \N__19114\,
            lcout => OPEN,
            ltout => \this_ppu.m9_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m9_0_a2_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19010\,
            in3 => \N__21242\,
            lcout => \this_ppu.N_97_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_0_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101011101010"
        )
    port map (
            in0 => \N__18980\,
            in1 => \N__19007\,
            in2 => \N__29791\,
            in3 => \N__28613\,
            lcout => \this_vga_signals.M_lcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_lcounter_q_RNI6R6E_0_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__18996\,
            in1 => \N__18978\,
            in2 => \_gnd_net_\,
            in3 => \N__35276\,
            lcout => \N_52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNI58DK1_5_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21164\,
            in1 => \N__20771\,
            in2 => \_gnd_net_\,
            in3 => \N__18968\,
            lcout => \this_ppu.N_814\,
            ltout => \this_ppu.N_814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIOVN89_10_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21341\,
            in2 => \N__18962\,
            in3 => \N__21949\,
            lcout => \this_ppu.N_806\,
            ltout => \this_ppu.N_806_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_2_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__30995\,
            in1 => \N__21435\,
            in2 => \N__18959\,
            in3 => \N__19124\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_5_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21438\,
            in1 => \N__19158\,
            in2 => \N__31018\,
            in3 => \N__19055\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_3_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19156\,
            in1 => \N__21436\,
            in2 => \N__31015\,
            in3 => \N__19103\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_4_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19157\,
            in1 => \N__21437\,
            in2 => \N__31016\,
            in3 => \N__19079\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_1_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__21434\,
            in1 => \N__19155\,
            in2 => \N__31017\,
            in3 => \N__19133\,
            lcout => \this_ppu.M_pixel_cnt_qZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21668\,
            in2 => \N__21235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21791\,
            in2 => \N__21278\,
            in3 => \N__19127\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_0\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_2_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21803\,
            in2 => \N__21296\,
            in3 => \N__19118\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_1\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_3_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19115\,
            in2 => \N__21908\,
            in3 => \N__19097\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_2\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19199\,
            in2 => \N__19094\,
            in3 => \N__19073\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_3\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_5_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19166\,
            in2 => \N__19070\,
            in3 => \N__19049\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_4\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_6_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21797\,
            in2 => \N__19046\,
            in3 => \N__19013\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_pixel_cnt_q_1_cry_5\,
            carryout => \this_ppu.un1_M_pixel_cnt_q_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_7_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__21991\,
            in1 => \N__21950\,
            in2 => \N__21262\,
            in3 => \N__19202\,
            lcout => \this_ppu.M_pixel_cnt_q_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_1_10_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21994\,
            in2 => \_gnd_net_\,
            in3 => \N__21947\,
            lcout => \this_ppu.M_state_q_RNISP3R6_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_10_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19193\,
            in2 => \_gnd_net_\,
            in3 => \N__23995\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_10_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__21948\,
            in1 => \_gnd_net_\,
            in2 => \N__21998\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_state_q_RNISP3R6Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_0_LC_12_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__23658\,
            in1 => \_gnd_net_\,
            in2 => \N__25198\,
            in3 => \N__23704\,
            lcout => \M_this_oam_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39391\,
            ce => 'H',
            sr => \N__38954\
        );

    \M_this_oam_address_q_3_LC_12_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__21898\,
            in1 => \N__19552\,
            in2 => \N__19594\,
            in3 => \N__25209\,
            lcout => \M_this_oam_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39395\,
            ce => 'H',
            sr => \N__38953\
        );

    \M_this_oam_address_q_4_LC_12_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19461\,
            in1 => \N__25200\,
            in2 => \_gnd_net_\,
            in3 => \N__19528\,
            lcout => \M_this_oam_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39395\,
            ce => 'H',
            sr => \N__38953\
        );

    \M_this_oam_address_q_5_LC_12_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__19529\,
            in1 => \N__19504\,
            in2 => \N__19468\,
            in3 => \N__25210\,
            lcout => \M_this_oam_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39395\,
            ce => 'H',
            sr => \N__38953\
        );

    \M_this_oam_address_q_2_LC_12_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__19551\,
            in1 => \N__25199\,
            in2 => \_gnd_net_\,
            in3 => \N__21897\,
            lcout => \M_this_oam_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39395\,
            ce => 'H',
            sr => \N__38953\
        );

    \M_this_oam_address_q_RNILNG41_3_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21899\,
            in1 => \N__19587\,
            in2 => \_gnd_net_\,
            in3 => \N__19550\,
            lcout => \un1_M_this_oam_address_q_c4\,
            ltout => \un1_M_this_oam_address_q_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIOKR51_5_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19503\,
            in2 => \N__19484\,
            in3 => \N__19460\,
            lcout => \un1_M_this_oam_address_q_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_0_1_LC_12_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__23758\,
            in1 => \N__23721\,
            in2 => \N__23671\,
            in3 => \N__36947\,
            lcout => \N_1240_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIMU531_LC_12_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23763\,
            in1 => \N__23662\,
            in2 => \_gnd_net_\,
            in3 => \N__23719\,
            lcout => \M_this_oam_ram_write_data_0_sqmuxa\,
            ltout => \M_this_oam_ram_write_data_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI32IG1_LC_12_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__37650\,
            in1 => \_gnd_net_\,
            in2 => \N__19409\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_write_data_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_LC_12_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__23764\,
            in1 => \N__23720\,
            in2 => \N__36965\,
            in3 => \N__23663\,
            lcout => \N_1232_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI4JDD1_LC_12_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19214\,
            in1 => \N__19266\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_oam_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_tmp_q_esr_0_LC_12_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38078\,
            lcout => \M_this_data_tmp_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39413\,
            ce => \N__23619\,
            sr => \N__36839\
        );

    \M_this_data_tmp_q_esr_4_LC_12_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37522\,
            lcout => \M_this_data_tmp_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39413\,
            ce => \N__23619\,
            sr => \N__36839\
        );

    \M_this_data_tmp_q_esr_2_LC_12_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37615\,
            lcout => \M_this_data_tmp_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39413\,
            ce => \N__23619\,
            sr => \N__36839\
        );

    \M_this_data_tmp_q_esr_21_LC_12_31_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38894\,
            lcout => \M_this_data_tmp_qZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39423\,
            ce => \N__21848\,
            sr => \N__36844\
        );

    \this_spr_ram.mem_mem_3_0_RNIQI5G_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19835\,
            in1 => \N__19811\,
            in2 => \_gnd_net_\,
            in3 => \N__20830\,
            lcout => \this_spr_ram.mem_mem_3_0_RNIQI5GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_0_0_RNIK6VF_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20824\,
            in1 => \N__19793\,
            in2 => \_gnd_net_\,
            in3 => \N__19778\,
            lcout => \this_spr_ram.mem_mem_0_0_RNIK6VFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_1_0_RNIMA1G_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19763\,
            in1 => \N__19742\,
            in2 => \_gnd_net_\,
            in3 => \N__20829\,
            lcout => \this_spr_ram.mem_mem_1_0_RNIMA1GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_RNIOE3G_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20828\,
            in1 => \N__19727\,
            in2 => \_gnd_net_\,
            in3 => \N__19709\,
            lcout => OPEN,
            ltout => \this_spr_ram.mem_mem_2_0_RNIOE3GZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIPCNI1_12_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__19692\,
            in1 => \N__19911\,
            in2 => \N__19655\,
            in3 => \N__19652\,
            lcout => \this_spr_ram.mem_DOUT_7_i_m2_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_RNIFL8S2_11_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__19646\,
            in1 => \N__19640\,
            in2 => \N__19928\,
            in3 => \N__19634\,
            lcout => \M_this_spr_ram_read_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_13_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20705\,
            in1 => \N__20690\,
            in2 => \_gnd_net_\,
            in3 => \N__32688\,
            lcout => \this_spr_ram.mem_radregZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI7SFJ1_3_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20681\,
            in1 => \N__20669\,
            in2 => \_gnd_net_\,
            in3 => \N__32664\,
            lcout => \M_this_ppu_spr_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI9TFJ1_4_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20441\,
            in1 => \N__20429\,
            in2 => \_gnd_net_\,
            in3 => \N__32663\,
            lcout => \M_this_ppu_spr_addr_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNIB6J72_8_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111000010100"
        )
    port map (
            in0 => \N__32665\,
            in1 => \N__24927\,
            in2 => \N__26567\,
            in3 => \N__24928\,
            lcout => \M_this_ppu_spr_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_1_RNIQE3G_0_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20838\,
            in1 => \N__19997\,
            in2 => \_gnd_net_\,
            in3 => \N__19982\,
            lcout => \this_spr_ram.mem_mem_2_1_RNIQE3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_radreg_11_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19961\,
            in1 => \N__19949\,
            in2 => \_gnd_net_\,
            in3 => \N__32669\,
            lcout => \this_spr_ram.mem_radregZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_4_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__22076\,
            in2 => \_gnd_net_\,
            in3 => \N__22151\,
            lcout => \this_ppu_M_screen_y_q_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39301\,
            ce => \N__23060\,
            sr => \N__36826\
        );

    \this_ppu.M_state_q_8_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000010001"
        )
    port map (
            in0 => \N__19856\,
            in1 => \N__36958\,
            in2 => \N__20741\,
            in3 => \N__20770\,
            lcout => \this_ppu.M_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39306\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m71_i_m2_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111011"
        )
    port map (
            in0 => \N__21375\,
            in1 => \N__21772\,
            in2 => \N__24049\,
            in3 => \N__20768\,
            lcout => \this_ppu.N_797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIFCA89_2_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23096\,
            in1 => \N__22119\,
            in2 => \_gnd_net_\,
            in3 => \N__22096\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c4\,
            ltout => \this_ppu.un3_M_screen_y_d_0_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIMH2E9_5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22385\,
            in2 => \N__20915\,
            in3 => \N__22085\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_4_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__30984\,
            in1 => \N__21099\,
            in2 => \N__20912\,
            in3 => \N__20996\,
            lcout => \this_ppu.M_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_1_RNISI5G_0_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20897\,
            in1 => \N__20882\,
            in2 => \_gnd_net_\,
            in3 => \N__20867\,
            lcout => \this_spr_ram.mem_mem_3_1_RNISI5GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_6_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20769\,
            in1 => \N__20737\,
            in2 => \_gnd_net_\,
            in3 => \N__36956\,
            lcout => \this_ppu.M_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_9_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__36955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20714\,
            lcout => \this_ppu.M_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39312\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNO_0_6_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__24164\,
            in2 => \N__21020\,
            in3 => \N__24305\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_surface_x_q_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_6_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__24086\,
            in1 => \N__22266\,
            in2 => \N__20708\,
            in3 => \N__21035\,
            lcout => \M_this_ppu_map_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39318\,
            ce => 'H',
            sr => \N__36819\
        );

    \this_ppu.M_state_q_ns_11_0__m35_i_o2_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__21170\,
            in1 => \N__21189\,
            in2 => \_gnd_net_\,
            in3 => \N__21091\,
            lcout => \this_ppu.N_798_0\,
            ltout => \this_ppu.N_798_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNIN4DCD_1_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__24574\,
            in1 => \N__24864\,
            in2 => \N__21023\,
            in3 => \N__24914\,
            lcout => \this_ppu.un1_M_surface_x_q_c3\,
            ltout => \this_ppu.un1_M_surface_x_q_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_3_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__21050\,
            in1 => \N__22267\,
            in2 => \N__21011\,
            in3 => \N__24306\,
            lcout => \M_this_ppu_map_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39318\,
            ce => 'H',
            sr => \N__36819\
        );

    \this_ppu.M_surface_x_q_0_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010011001"
        )
    port map (
            in0 => \N__24915\,
            in1 => \N__21008\,
            in2 => \N__21398\,
            in3 => \N__22268\,
            lcout => \this_ppu.offset_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39318\,
            ce => 'H',
            sr => \N__36819\
        );

    \this_ppu.M_surface_x_q_RNO_0_7_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22285\,
            in1 => \N__24163\,
            in2 => \N__24093\,
            in3 => \N__24243\,
            lcout => \this_ppu.un1_M_surface_x_q_ac0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNINHSUC_1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__24863\,
            in1 => \N__20992\,
            in2 => \N__21116\,
            in3 => \N__24913\,
            lcout => \this_ppu.un1_M_surface_x_q_c2\,
            ltout => \this_ppu.un1_M_surface_x_q_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNO_0_5_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24304\,
            in1 => \N__24245\,
            in2 => \N__21002\,
            in3 => \N__24572\,
            lcout => OPEN,
            ltout => \this_ppu.un1_M_surface_x_q_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_5_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__21041\,
            in1 => \N__22252\,
            in2 => \N__20999\,
            in3 => \N__24165\,
            lcout => \M_this_ppu_map_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39326\,
            ce => 'H',
            sr => \N__36816\
        );

    \this_ppu.M_state_q_RNII1FQB_7_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__21155\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21190\,
            lcout => \this_ppu.N_800\,
            ltout => \this_ppu.N_800_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNICH7OC_11_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21112\,
            in1 => \N__26690\,
            in2 => \N__20981\,
            in3 => \N__20975\,
            lcout => \N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_2_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22251\,
            in1 => \N__21197\,
            in2 => \N__21062\,
            in3 => \N__24573\,
            lcout => \this_ppu.M_surface_x_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39326\,
            ce => 'H',
            sr => \N__36816\
        );

    \this_ppu.M_state_q_RNIOVBHC_7_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__21191\,
            in1 => \N__21156\,
            in2 => \N__21115\,
            in3 => \N__24912\,
            lcout => \this_ppu.un1_M_surface_x_q_c1\,
            ltout => \this_ppu.un1_M_surface_x_q_c1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_RNIOOTPD_1_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24303\,
            in1 => \N__24571\,
            in2 => \N__21065\,
            in3 => \N__24862\,
            lcout => \this_ppu.un1_M_surface_x_q_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_10_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37652\,
            lcout => \M_this_scroll_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_11_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37898\,
            lcout => \M_this_scroll_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_12_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_13_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38910\,
            lcout => \M_this_scroll_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_14_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_15_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38760\,
            lcout => \M_this_scroll_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_8_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38129\,
            lcout => \M_this_scroll_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \M_this_scroll_q_esr_9_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37739\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39334\,
            ce => \N__23501\,
            sr => \N__36820\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIFICF2_5_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__33172\,
            in1 => \N__23531\,
            in2 => \_gnd_net_\,
            in3 => \N__33942\,
            lcout => OPEN,
            ltout => \N_829_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m14_0_o2_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000001"
        )
    port map (
            in0 => \N__34073\,
            in1 => \N__34650\,
            in2 => \N__21383\,
            in3 => \N__34752\,
            lcout => \N_58_0\,
            ltout => \N_58_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI4GQN4_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__29810\,
            in1 => \N__21594\,
            in2 => \N__21380\,
            in3 => \N__29847\,
            lcout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0\,
            ltout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_7_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__21643\,
            in1 => \N__21372\,
            in2 => \N__21305\,
            in3 => \N__21302\,
            lcout => \this_ppu.M_pixel_cnt_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39342\,
            ce => 'H',
            sr => \N__36822\
        );

    \this_ppu.M_state_q_ns_11_0__m9_0_a2_4_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21295\,
            in1 => \N__21274\,
            in2 => \N__21263\,
            in3 => \N__21231\,
            lcout => \this_ppu.m9_0_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_pixel_cnt_q_RNO_0_0_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__21980\,
            in1 => \N__21236\,
            in2 => \_gnd_net_\,
            in3 => \N__21945\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNIJ1SE_10_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__21710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21777\,
            lcout => \this_ppu.N_60_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_2_10_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21943\,
            lcout => \this_ppu.M_state_q_RNISP3R6_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_4_10_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21944\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21979\,
            lcout => \this_ppu.M_state_q_RNISP3R6_4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_0_10_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21942\,
            lcout => \this_ppu.M_state_q_RNISP3R6_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_RNI5CEE4_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__29809\,
            in1 => \N__29848\,
            in2 => \_gnd_net_\,
            in3 => \N__29821\,
            lcout => \this_ppu.N_835_0\,
            ltout => \this_ppu.N_835_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNINHM65_10_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__21709\,
            in2 => \N__21674\,
            in3 => \N__21608\,
            lcout => \this_ppu.N_783\,
            ltout => \this_ppu.N_783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNO_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21671\,
            in3 => \N__21976\,
            lcout => \this_ppu.un1_M_pixel_cnt_q_1_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIDQQ11_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36546\,
            in2 => \_gnd_net_\,
            in3 => \N__36170\,
            lcout => \N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_2_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21662\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39360\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_0_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21993\,
            in1 => \N__21639\,
            in2 => \N__21621\,
            in3 => \N__21476\,
            lcout => \this_ppu.N_807\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_RNISP3R6_3_10_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21992\,
            in2 => \_gnd_net_\,
            in3 => \N__21946\,
            lcout => \this_ppu.M_state_q_RNISP3R6_3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIR9R11_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__25943\,
            in1 => \N__25253\,
            in2 => \N__25304\,
            in3 => \N__34931\,
            lcout => \N_222_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNIMU531_1_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23693\,
            in1 => \N__36545\,
            in2 => \N__23765\,
            in3 => \N__34926\,
            lcout => \un1_M_this_oam_address_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_1_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__23667\,
            in1 => \N__23759\,
            in2 => \N__25216\,
            in3 => \N__23723\,
            lcout => \M_this_oam_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39396\,
            ce => 'H',
            sr => \N__38951\
        );

    \M_this_data_tmp_q_esr_18_LC_13_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39402\,
            ce => \N__21825\,
            sr => \N__36834\
        );

    \M_this_data_tmp_q_esr_1_LC_13_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_tmp_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39409\,
            ce => \N__23606\,
            sr => \N__36836\
        );

    \M_this_data_tmp_q_esr_19_LC_13_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37852\,
            lcout => \M_this_data_tmp_qZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39417\,
            ce => \N__21849\,
            sr => \N__36840\
        );

    \this_ppu.M_screen_y_q_esr_3_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__23094\,
            in1 => \N__22097\,
            in2 => \N__22134\,
            in3 => \N__23178\,
            lcout => \this_ppu_M_screen_y_q_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39302\,
            ce => \N__23059\,
            sr => \N__36823\
        );

    \this_ppu.M_screen_y_q_esr_6_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22355\,
            in1 => \N__22162\,
            in2 => \_gnd_net_\,
            in3 => \N__23180\,
            lcout => \this_ppu_M_screen_y_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39302\,
            ce => \N__23059\,
            sr => \N__36823\
        );

    \this_ppu.M_screen_y_q_esr_7_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100010100000"
        )
    port map (
            in0 => \N__23181\,
            in1 => \N__22356\,
            in2 => \N__23320\,
            in3 => \N__22163\,
            lcout => \this_ppu.M_screen_y_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39302\,
            ce => \N__23059\,
            sr => \N__36823\
        );

    \this_ppu.M_screen_y_q_esr_5_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__22077\,
            in1 => \N__22150\,
            in2 => \N__22396\,
            in3 => \N__23179\,
            lcout => \this_ppu_M_screen_y_q_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39302\,
            ce => \N__23059\,
            sr => \N__36823\
        );

    \this_ppu.M_screen_y_q_esr_RNIO9AV8_3_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__23140\,
            in1 => \N__22118\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIO9AV8Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_RNICCMV8_0_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23254\,
            in2 => \_gnd_net_\,
            in3 => \N__23139\,
            lcout => \this_ppu.M_screen_y_q_RNICCMV8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNICBI29_1_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23209\,
            in1 => \N__23253\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \this_ppu.un3_M_screen_y_d_0_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIN8AV8_2_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23090\,
            in2 => \_gnd_net_\,
            in3 => \N__23141\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIN8AV8Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIPAAV8_4_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23142\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22084\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIPAAV8Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m68_0_a2_2_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__22043\,
            in1 => \N__24275\,
            in2 => \_gnd_net_\,
            in3 => \N__24059\,
            lcout => OPEN,
            ltout => \this_ppu.m68_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_state_q_ns_11_0__m68_0_a2_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24209\,
            in1 => \N__24131\,
            in2 => \N__22022\,
            in3 => \N__25010\,
            lcout => \this_ppu.M_state_q_ns_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIM8ES8_9_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34153\,
            in2 => \_gnd_net_\,
            in3 => \N__29607\,
            lcout => \M_this_ppu_vga_is_drawing\,
            ltout => \M_this_ppu_vga_is_drawing_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIM7AV8_1_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22400\,
            in3 => \N__23210\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIM7AV8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIQBAV8_5_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23143\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIQBAV8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_esr_RNIRCAV8_6_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22357\,
            lcout => \this_ppu.M_screen_y_q_esr_RNIRCAV8Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_x_q_1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__22334\,
            in1 => \N__22255\,
            in2 => \N__22328\,
            in3 => \N__24865\,
            lcout => \this_ppu.M_surface_x_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39319\,
            ce => 'H',
            sr => \N__36813\
        );

    \this_ppu.line_clk.M_last_q_RNIGL6V4_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__22253\,
            in1 => \_gnd_net_\,
            in2 => \N__36964\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.M_oam_cache_cnt_d_0_sqmuxa_i_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_screen_y_q_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__23158\,
            in1 => \N__23241\,
            in2 => \N__23257\,
            in3 => \N__22257\,
            lcout => \M_this_ppu_vram_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39319\,
            ce => 'H',
            sr => \N__36813\
        );

    \this_ppu.M_surface_x_q_7_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__22254\,
            in1 => \N__25045\,
            in2 => \N__22313\,
            in3 => \N__22304\,
            lcout => \M_this_ppu_map_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39319\,
            ce => 'H',
            sr => \N__36813\
        );

    \this_ppu.M_surface_x_q_4_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__22295\,
            in1 => \N__22286\,
            in2 => \N__24253\,
            in3 => \N__22256\,
            lcout => \M_this_ppu_map_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39319\,
            ce => 'H',
            sr => \N__36813\
        );

    \this_ppu.oam_cache.read_data_RNI6RFJ1_2_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22190\,
            in1 => \N__22178\,
            in2 => \_gnd_net_\,
            in3 => \N__32687\,
            lcout => \M_this_ppu_spr_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CRY_0_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23171\,
            in2 => \N__23183\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.M_surface_y_q_esr_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22751\,
            in2 => \N__25004\,
            in3 => \N__22706\,
            lcout => \this_ppu.offset_y\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_0_0_c_THRU_CO\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_0\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_1_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22703\,
            in2 => \N__24995\,
            in3 => \N__22667\,
            lcout => \this_ppu.M_surface_y_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_0\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_1\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_2_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22664\,
            in2 => \N__24986\,
            in3 => \N__22625\,
            lcout => \this_ppu.M_surface_y_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_1\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_2\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_3_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22622\,
            in2 => \N__24977\,
            in3 => \N__22568\,
            lcout => \M_this_ppu_map_addr_5\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_2\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_3\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_4_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22565\,
            in2 => \N__24965\,
            in3 => \N__22517\,
            lcout => \M_this_ppu_map_addr_6\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_3\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_4\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_5_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22514\,
            in2 => \N__24956\,
            in3 => \N__22457\,
            lcout => \M_this_ppu_map_addr_7\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_4\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_5\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_6_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22454\,
            in2 => \N__24947\,
            in3 => \N__23327\,
            lcout => \M_this_ppu_map_addr_8\,
            ltout => OPEN,
            carryin => \this_ppu.un1_M_surface_y_d_cry_5\,
            carryout => \this_ppu.un1_M_surface_y_d_cry_6\,
            clk => \N__39327\,
            ce => \N__23058\,
            sr => \N__36817\
        );

    \this_ppu.M_surface_y_q_esr_7_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__23177\,
            in1 => \N__24938\,
            in2 => \N__23324\,
            in3 => \N__23303\,
            lcout => \M_this_ppu_map_addr_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39335\,
            ce => \N__23051\,
            sr => \N__36821\
        );

    \this_ppu.M_screen_y_q_esr_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__23255\,
            in1 => \N__23207\,
            in2 => \_gnd_net_\,
            in3 => \N__23175\,
            lcout => \this_ppu.M_screen_y_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39335\,
            ce => \N__23051\,
            sr => \N__36821\
        );

    \this_ppu.M_screen_y_q_esr_2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100000000000"
        )
    port map (
            in0 => \N__23256\,
            in1 => \N__23208\,
            in2 => \N__23095\,
            in3 => \N__23176\,
            lcout => \this_ppu.M_screen_y_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39335\,
            ce => \N__23051\,
            sr => \N__36821\
        );

    \CONSTANT_ONE_LUT4_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIP7R11_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__25941\,
            in1 => \N__25248\,
            in2 => \N__25300\,
            in3 => \N__34994\,
            lcout => \M_this_state_d_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25291\,
            lcout => \this_start_data_delay.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__25292\,
            in1 => \N__25937\,
            in2 => \_gnd_net_\,
            in3 => \N__25247\,
            lcout => \this_start_data_delay.N_227_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_11_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23021\,
            in2 => \_gnd_net_\,
            in3 => \N__24001\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_delay_clk.M_pipe_q_4_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23519\,
            lcout => \M_this_delay_clk_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNILR691_2_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__36498\,
            in1 => \N__36943\,
            in2 => \_gnd_net_\,
            in3 => \N__36065\,
            lcout => \N_1256_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_1_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__25130\,
            in1 => \N__26759\,
            in2 => \_gnd_net_\,
            in3 => \N__25882\,
            lcout => \M_this_data_count_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39353\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_2_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__26760\,
            in1 => \N__25115\,
            in2 => \_gnd_net_\,
            in3 => \N__25903\,
            lcout => \M_this_data_count_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39353\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_3_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__25103\,
            in1 => \N__26761\,
            in2 => \_gnd_net_\,
            in3 => \N__25860\,
            lcout => \M_this_data_count_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39353\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_7_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__26762\,
            in1 => \_gnd_net_\,
            in2 => \N__25082\,
            in3 => \N__26880\,
            lcout => \M_this_data_count_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39353\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23997\,
            in2 => \_gnd_net_\,
            in3 => \N__23489\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_0_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23998\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23444\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_1_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23999\,
            in2 => \_gnd_net_\,
            in3 => \N__23402\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.mem_mem_0_1_RNO_10_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24000\,
            in1 => \N__23354\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ctrl_flags_q_6_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24036\,
            in1 => \N__36544\,
            in2 => \N__37375\,
            in3 => \N__36032\,
            lcout => \M_this_ctrl_flags_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39361\,
            ce => 'H',
            sr => \N__36827\
        );

    \this_ppu.oam_cache.mem_mem_0_0_RNO_12_LC_14_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24017\,
            in2 => \_gnd_net_\,
            in3 => \N__23996\,
            lcout => \this_ppu.oam_cache.M_oam_cache_write_data_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_oam_address_q_RNI24IA1_1_1_LC_14_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__23757\,
            in1 => \N__23722\,
            in2 => \N__23672\,
            in3 => \N__36934\,
            lcout => \N_1248_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_2_LC_14_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25820\,
            lcout => \this_reset_cond.M_stage_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_3_LC_14_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30818\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23573\,
            lcout => \this_reset_cond.M_stage_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK6R81_1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__36539\,
            in1 => \N__35633\,
            in2 => \_gnd_net_\,
            in3 => \N__38277\,
            lcout => \M_this_spr_ram_write_en_0_i_1_0\,
            ltout => \M_this_spr_ram_write_en_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_6_0_wclke_3_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32000\,
            in1 => \N__32204\,
            in2 => \N__23567\,
            in3 => \N__32102\,
            lcout => \this_spr_ram.mem_WE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIQVHO1_0_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__31226\,
            in1 => \N__26535\,
            in2 => \N__31354\,
            in3 => \N__26659\,
            lcout => \this_vga_signals.M_vcounter_d7lt8_0\,
            ltout => \this_vga_signals.M_vcounter_d7lt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI542T3_9_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__26393\,
            in1 => \N__33940\,
            in2 => \N__24932\,
            in3 => \N__35271\,
            lcout => \this_vga_signals.M_vcounter_d8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_0_c_inv_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24884\,
            in2 => \N__24929\,
            in3 => \N__26554\,
            lcout => \this_ppu.M_oam_cache_read_data_i_8\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \this_ppu.offset_x_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_0_c_RNI5N4U1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__32680\,
            in1 => \N__24878\,
            in2 => \N__24866\,
            in3 => \N__24590\,
            lcout => \M_this_ppu_spr_addr_1\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_0\,
            carryout => \this_ppu.offset_x_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_1_c_RNIFSQU1_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__32694\,
            in1 => \N__24587\,
            in2 => \N__24578\,
            in3 => \N__24332\,
            lcout => \M_this_ppu_spr_addr_2\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_1\,
            carryout => \this_ppu.offset_x_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_2_c_RNI0QAP_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26363\,
            in2 => \N__24328\,
            in3 => \N__24269\,
            lcout => \this_ppu.offset_x_3\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_2\,
            carryout => \this_ppu.offset_x_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_3_c_RNI3UBP_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26591\,
            in2 => \N__24252\,
            in3 => \N__24203\,
            lcout => \this_ppu.offset_x_4\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_3\,
            carryout => \this_ppu.offset_x_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_4_c_RNI62DP_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24200\,
            in2 => \N__24181\,
            in3 => \N__24125\,
            lcout => \this_ppu.offset_x_5\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_4\,
            carryout => \this_ppu.offset_x_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_5_c_RNI96EP_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24122\,
            in2 => \N__24103\,
            in3 => \N__24053\,
            lcout => \this_ppu.offset_x_6\,
            ltout => OPEN,
            carryin => \this_ppu.offset_x_cry_5\,
            carryout => \this_ppu.offset_x_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.offset_x_cry_6_c_RNICAFP_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__25044\,
            in1 => \_gnd_net_\,
            in2 => \N__25025\,
            in3 => \N__25013\,
            lcout => \this_ppu.offset_x_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_scroll_q_esr_0_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38128\,
            lcout => \M_this_scroll_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_1_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37759\,
            lcout => \M_this_scroll_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_2_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37628\,
            lcout => \M_this_scroll_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_3_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37879\,
            lcout => \M_this_scroll_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_4_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_5_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38890\,
            lcout => \M_this_scroll_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_6_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37351\,
            lcout => \M_this_scroll_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_scroll_q_esr_7_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__38759\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \M_this_scroll_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39320\,
            ce => \N__35522\,
            sr => \N__36814\
        );

    \M_this_data_count_q_cry_c_0_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25838\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_19_0_\,
            carryout => \M_this_data_count_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_0_THRU_LUT4_0_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25883\,
            in2 => \N__25402\,
            in3 => \N__25118\,
            lcout => \M_this_data_count_q_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_0\,
            carryout => \M_this_data_count_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_1_THRU_LUT4_0_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25370\,
            in2 => \N__25907\,
            in3 => \N__25106\,
            lcout => \M_this_data_count_q_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_1\,
            carryout => \M_this_data_count_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_2_THRU_LUT4_0_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25862\,
            in2 => \N__25403\,
            in3 => \N__25094\,
            lcout => \M_this_data_count_q_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_2\,
            carryout => \M_this_data_count_q_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_3_THRU_LUT4_0_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25374\,
            in2 => \N__26021\,
            in3 => \N__25091\,
            lcout => \M_this_data_count_q_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_3\,
            carryout => \M_this_data_count_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_4_THRU_LUT4_0_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25988\,
            in2 => \N__25404\,
            in3 => \N__25088\,
            lcout => \M_this_data_count_q_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_4\,
            carryout => \M_this_data_count_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_5_THRU_LUT4_0_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25378\,
            in2 => \N__26714\,
            in3 => \N__25085\,
            lcout => \M_this_data_count_q_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_5\,
            carryout => \M_this_data_count_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_6_THRU_LUT4_0_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26882\,
            in2 => \N__25405\,
            in3 => \N__25070\,
            lcout => \M_this_data_count_q_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_6\,
            carryout => \M_this_data_count_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_8_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25142\,
            in2 => \N__25400\,
            in3 => \N__25067\,
            lcout => \M_this_data_count_q_s_8\,
            ltout => OPEN,
            carryin => \bfn_15_20_0_\,
            carryout => \M_this_data_count_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_8_THRU_LUT4_0_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25366\,
            in2 => \N__25964\,
            in3 => \N__25814\,
            lcout => \M_this_data_count_q_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_8\,
            carryout => \M_this_data_count_q_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_10_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26792\,
            in2 => \N__25399\,
            in3 => \N__25811\,
            lcout => \M_this_data_count_q_s_10\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_9\,
            carryout => \M_this_data_count_q_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_10_THRU_LUT4_0_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25362\,
            in2 => \N__26825\,
            in3 => \N__25808\,
            lcout => \M_this_data_count_q_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_10\,
            carryout => \M_this_data_count_q_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_cry_11_THRU_LUT4_0_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26840\,
            in2 => \N__25401\,
            in3 => \N__25310\,
            lcout => \M_this_data_count_q_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \M_this_data_count_q_cry_11\,
            carryout => \M_this_data_count_q_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_RNO_0_13_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26806\,
            in2 => \_gnd_net_\,
            in3 => \N__25307\,
            lcout => \M_this_data_count_q_s_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBJQQ_0_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__25296\,
            in1 => \N__25936\,
            in2 => \_gnd_net_\,
            in3 => \N__25246\,
            lcout => \N_220_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_9_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36502\,
            in1 => \N__36957\,
            in2 => \_gnd_net_\,
            in3 => \N__35621\,
            lcout => \M_this_state_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_8_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__36949\,
            in1 => \N__25226\,
            in2 => \N__25211\,
            in3 => \N__26753\,
            lcout => \M_this_data_count_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39344\,
            ce => \N__32294\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_7_11_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25141\,
            in1 => \N__25983\,
            in2 => \N__25963\,
            in3 => \N__26013\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_a2_0_7Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_4_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__26014\,
            in1 => \N__26033\,
            in2 => \_gnd_net_\,
            in3 => \N__26750\,
            lcout => \M_this_data_count_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39344\,
            ce => \N__32294\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_5_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000101"
        )
    port map (
            in0 => \N__26751\,
            in1 => \_gnd_net_\,
            in2 => \N__26000\,
            in3 => \N__25984\,
            lcout => \M_this_data_count_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39344\,
            ce => \N__32294\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_9_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__25970\,
            in1 => \N__26752\,
            in2 => \_gnd_net_\,
            in3 => \N__25959\,
            lcout => \M_this_data_count_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39344\,
            ce => \N__32294\,
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI30CP2_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__38308\,
            in1 => \N__25942\,
            in2 => \_gnd_net_\,
            in3 => \N__36948\,
            lcout => \N_685_i\,
            ltout => \N_685_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_0_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001001"
        )
    port map (
            in0 => \N__25834\,
            in1 => \_gnd_net_\,
            in2 => \N__25910\,
            in3 => \_gnd_net_\,
            lcout => \M_this_data_count_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39344\,
            ce => \N__32294\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_9_11_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25899\,
            in1 => \N__25878\,
            in2 => \N__25861\,
            in3 => \N__25833\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_a2_0_9Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_5_LC_15_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26336\,
            in2 => \_gnd_net_\,
            in3 => \N__30801\,
            lcout => \this_reset_cond.M_stage_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_1_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30815\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26330\,
            lcout => \this_reset_cond.M_stage_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_4_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30816\,
            in2 => \_gnd_net_\,
            in3 => \N__26342\,
            lcout => \this_reset_cond.M_stage_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_0_LC_15_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_reset_cond.M_stage_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI4PFJ1_0_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26051\,
            in1 => \N__26324\,
            in2 => \_gnd_net_\,
            in3 => \N__32701\,
            lcout => \M_this_ppu_spr_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_0_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26066\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39288\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29770\,
            in1 => \N__26536\,
            in2 => \N__28616\,
            in3 => \N__28611\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            clk => \N__39296\,
            ce => 'H',
            sr => \N__34426\
        );

    \this_vga_signals.M_vcounter_q_1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29772\,
            in1 => \N__26666\,
            in2 => \_gnd_net_\,
            in3 => \N__26045\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_0\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            clk => \N__39296\,
            ce => 'H',
            sr => \N__34426\
        );

    \this_vga_signals.M_vcounter_q_2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29771\,
            in1 => \N__31260\,
            in2 => \_gnd_net_\,
            in3 => \N__26042\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_1\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            clk => \N__39296\,
            ce => 'H',
            sr => \N__34426\
        );

    \this_vga_signals.M_vcounter_q_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__29773\,
            in1 => \N__31352\,
            in2 => \_gnd_net_\,
            in3 => \N__26039\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_3\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_2\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            clk => \N__39296\,
            ce => 'H',
            sr => \N__34426\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OH_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33941\,
            in2 => \_gnd_net_\,
            in3 => \N__26036\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_3_c_RNIJ5OHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_3\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PH_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33184\,
            in2 => \_gnd_net_\,
            in3 => \N__26408\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_4_c_RNIL8PHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_4\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQH_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34061\,
            in2 => \_gnd_net_\,
            in3 => \N__26405\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_5_c_RNINBQHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_5\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERH_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34754\,
            in2 => \_gnd_net_\,
            in3 => \N__26402\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_6_c_RNIPERHZ0\,
            ltout => OPEN,
            carryin => \this_vga_signals.un1_M_vcounter_q_cry_6\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSH_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34655\,
            in3 => \N__26399\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_7_c_RNIRHSHZ0\,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \this_vga_signals.un1_M_vcounter_q_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTH_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35272\,
            in2 => \_gnd_net_\,
            in3 => \N__26396\,
            lcout => \this_vga_signals.un1_M_vcounter_q_cry_8_c_RNITKTHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNILL3J1_1_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31353\,
            in1 => \N__26667\,
            in2 => \N__34753\,
            in3 => \N__33925\,
            lcout => \this_vga_signals.m43_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIIDLD1_7_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34060\,
            in1 => \N__34651\,
            in2 => \N__33183\,
            in3 => \N__34745\,
            lcout => \this_vga_signals.M_vcounter_d7lto9_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIPIAB9_9_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__28538\,
            in1 => \N__34154\,
            in2 => \_gnd_net_\,
            in3 => \N__29598\,
            lcout => port_nmib_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI72M7_11_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26609\,
            lcout => \this_ppu.M_oam_cache_read_data_i_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_11_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26357\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39305\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI83M7_12_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26603\,
            lcout => \this_ppu.M_oam_cache_read_data_i_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_8_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26585\,
            lcout => \this_ppu.M_oam_cache_read_data_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_N_2L1_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000100"
        )
    port map (
            in0 => \N__30488\,
            in1 => \N__31523\,
            in2 => \_gnd_net_\,
            in3 => \N__30581\,
            lcout => \this_vga_signals.g0_41_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100001000111"
        )
    port map (
            in0 => \N__30417\,
            in1 => \N__29966\,
            in2 => \N__30287\,
            in3 => \N__26504\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_15_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010110000101"
        )
    port map (
            in0 => \N__26669\,
            in1 => \N__26543\,
            in2 => \N__26519\,
            in3 => \N__31187\,
            lcout => \this_vga_signals.mult1_un82_sum_c3_0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_N_4L5_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010101111"
        )
    port map (
            in0 => \N__31405\,
            in1 => \_gnd_net_\,
            in2 => \N__30419\,
            in3 => \N__30002\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_41_N_4L5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_1_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31286\,
            in1 => \N__26516\,
            in2 => \N__26507\,
            in3 => \N__29891\,
            lcout => \this_vga_signals.g0_41_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNI8D7RUG1_2_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__30047\,
            in1 => \N__29912\,
            in2 => \N__26498\,
            in3 => \N__26432\,
            lcout => \M_this_vga_signals_address_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIVIOMG4_2_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000111011"
        )
    port map (
            in0 => \N__31287\,
            in1 => \N__29996\,
            in2 => \N__26624\,
            in3 => \N__31406\,
            lcout => \this_vga_signals.mult1_un68_sum_c3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x2_4_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30501\,
            in1 => \N__30223\,
            in2 => \N__30017\,
            in3 => \N__30590\,
            lcout => \this_vga_signals.g0_i_x2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__31739\,
            in1 => \N__31094\,
            in2 => \N__30230\,
            in3 => \N__29960\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_c3_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101110111101"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__31288\,
            in2 => \N__26636\,
            in3 => \N__26633\,
            lcout => \this_vga_signals.if_m5_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBOQ11_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38171\,
            lcout => \N_241_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_18_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000010"
        )
    port map (
            in0 => \N__33608\,
            in1 => \N__33410\,
            in2 => \N__33185\,
            in3 => \N__30623\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_3_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__33938\,
            in1 => \_gnd_net_\,
            in2 => \N__26627\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI2UNG73_4_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101100101"
        )
    port map (
            in0 => \N__29906\,
            in1 => \N__31738\,
            in2 => \N__33209\,
            in3 => \N__30222\,
            lcout => \this_vga_signals.N_17_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g2_1_2_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__33409\,
            in1 => \N__34045\,
            in2 => \N__33944\,
            in3 => \N__33607\,
            lcout => \this_vga_signals.g2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_10_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__26757\,
            in1 => \N__26615\,
            in2 => \N__39530\,
            in3 => \N__36961\,
            lcout => \M_this_data_count_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39330\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_12_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__26900\,
            in1 => \N__26755\,
            in2 => \_gnd_net_\,
            in3 => \N__26839\,
            lcout => \M_this_data_count_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39330\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_13_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__26758\,
            in1 => \N__26894\,
            in2 => \N__35777\,
            in3 => \N__36962\,
            lcout => \M_this_data_count_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39330\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_11_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__26821\,
            in1 => \N__26888\,
            in2 => \_gnd_net_\,
            in3 => \N__26754\,
            lcout => \M_this_data_count_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39330\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_6_11_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26881\,
            in2 => \_gnd_net_\,
            in3 => \N__26703\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_this_state_q_srsts_i_a2_0_6Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_11_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26858\,
            in1 => \N__26780\,
            in2 => \N__26849\,
            in3 => \N__26846\,
            lcout => \N_930\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_q_srsts_i_a2_0_8_11_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26838\,
            in1 => \N__26820\,
            in2 => \N__26807\,
            in3 => \N__26791\,
            lcout => \this_vga_signals.M_this_state_q_srsts_i_a2_0_8Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_data_count_q_6_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__26704\,
            in1 => \_gnd_net_\,
            in2 => \N__26774\,
            in3 => \N__26756\,
            lcout => \M_this_data_count_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39330\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \M_this_ctrl_flags_q_5_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__26683\,
            in1 => \N__36551\,
            in2 => \N__38909\,
            in3 => \N__36034\,
            lcout => \M_this_ctrl_flags_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39338\,
            ce => 'H',
            sr => \N__36824\
        );

    \M_this_ctrl_flags_q_7_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__36033\,
            in1 => \N__38761\,
            in2 => \N__28534\,
            in3 => \N__36552\,
            lcout => \M_this_ctrl_flags_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39338\,
            ce => 'H',
            sr => \N__36824\
        );

    \this_reset_cond.M_stage_q_6_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28517\,
            lcout => \this_reset_cond.M_stage_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_spr_address_q_0_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35806\,
            in1 => \N__28302\,
            in2 => \N__28673\,
            in3 => \N__28672\,
            lcout => \M_this_spr_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \un1_M_this_spr_address_q_cry_0\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_1_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35810\,
            in1 => \N__28073\,
            in2 => \_gnd_net_\,
            in3 => \N__28058\,
            lcout => \M_this_spr_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_0\,
            carryout => \un1_M_this_spr_address_q_cry_1\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_2_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35807\,
            in1 => \N__27859\,
            in2 => \_gnd_net_\,
            in3 => \N__27809\,
            lcout => \M_this_spr_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_1\,
            carryout => \un1_M_this_spr_address_q_cry_2\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_3_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35811\,
            in1 => \N__27600\,
            in2 => \_gnd_net_\,
            in3 => \N__27569\,
            lcout => \M_this_spr_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_2\,
            carryout => \un1_M_this_spr_address_q_cry_3\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_4_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35808\,
            in1 => \N__27371\,
            in2 => \_gnd_net_\,
            in3 => \N__27347\,
            lcout => \M_this_spr_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_3\,
            carryout => \un1_M_this_spr_address_q_cry_4\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_5_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35812\,
            in1 => \N__27182\,
            in2 => \_gnd_net_\,
            in3 => \N__27140\,
            lcout => \M_this_spr_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_4\,
            carryout => \un1_M_this_spr_address_q_cry_5\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_6_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35809\,
            in1 => \N__26928\,
            in2 => \_gnd_net_\,
            in3 => \N__26903\,
            lcout => \M_this_spr_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_5\,
            carryout => \un1_M_this_spr_address_q_cry_6\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_7_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35813\,
            in1 => \N__29401\,
            in2 => \_gnd_net_\,
            in3 => \N__29357\,
            lcout => \M_this_spr_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_6\,
            carryout => \un1_M_this_spr_address_q_cry_7\,
            clk => \N__39290\,
            ce => 'H',
            sr => \N__38961\
        );

    \M_this_spr_address_q_8_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35783\,
            in1 => \N__29192\,
            in2 => \_gnd_net_\,
            in3 => \N__29150\,
            lcout => \M_this_spr_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_13_0_\,
            carryout => \un1_M_this_spr_address_q_cry_8\,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \M_this_spr_address_q_9_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35786\,
            in1 => \N__28959\,
            in2 => \_gnd_net_\,
            in3 => \N__28916\,
            lcout => \M_this_spr_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_8\,
            carryout => \un1_M_this_spr_address_q_cry_9\,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \M_this_spr_address_q_10_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35781\,
            in1 => \N__28722\,
            in2 => \_gnd_net_\,
            in3 => \N__28685\,
            lcout => \M_this_spr_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_9\,
            carryout => \un1_M_this_spr_address_q_cry_10\,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \M_this_spr_address_q_11_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35785\,
            in1 => \N__32080\,
            in2 => \_gnd_net_\,
            in3 => \N__28682\,
            lcout => \M_this_spr_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_10\,
            carryout => \un1_M_this_spr_address_q_cry_11\,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \M_this_spr_address_q_12_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35782\,
            in1 => \N__32176\,
            in2 => \_gnd_net_\,
            in3 => \N__28679\,
            lcout => \M_this_spr_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_spr_address_q_cry_11\,
            carryout => \un1_M_this_spr_address_q_cry_12\,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \M_this_spr_address_q_13_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31972\,
            in1 => \N__35784\,
            in2 => \_gnd_net_\,
            in3 => \N__28676\,
            lcout => \M_this_spr_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39293\,
            ce => 'H',
            sr => \N__38958\
        );

    \this_start_data_delay.M_last_q_RNIK6R81_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__38282\,
            in1 => \N__36567\,
            in2 => \_gnd_net_\,
            in3 => \N__35629\,
            lcout => \M_this_spr_ram_write_en_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNINK957_9_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28647\,
            in1 => \N__28610\,
            in2 => \_gnd_net_\,
            in3 => \N__29766\,
            lcout => \this_vga_signals.M_vcounter_q_esr_RNINK957Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIOLTE3_2_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__29885\,
            in1 => \N__30086\,
            in2 => \N__31272\,
            in3 => \N__34041\,
            lcout => this_vga_signals_vsync_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.line_clk.M_last_q_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29855\,
            in2 => \_gnd_net_\,
            in3 => \N__29828\,
            lcout => \this_ppu.line_clk.M_last_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39307\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNICF6E7_9_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29790\,
            in2 => \_gnd_net_\,
            in3 => \N__29650\,
            lcout => \this_vga_signals.N_933_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_36_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__33123\,
            in1 => \N__33000\,
            in2 => \_gnd_net_\,
            in3 => \N__32935\,
            lcout => \this_vga_signals.N_10_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_1_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_ppu.oam_cache.M_oam_cache_read_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39313\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIB4G42_9_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__34633\,
            in1 => \N__35257\,
            in2 => \N__30080\,
            in3 => \N__34732\,
            lcout => OPEN,
            ltout => \this_vga_signals.vvisibility_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIEK4D3_9_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29621\,
            in3 => \N__31159\,
            lcout => \this_vga_signals.vvisibility\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_4_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33687\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39321\,
            ce => \N__34484\,
            sr => \N__34427\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_0_1_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001011111"
        )
    port map (
            in0 => \N__33907\,
            in1 => \N__33126\,
            in2 => \N__34065\,
            in3 => \N__33610\,
            lcout => \this_vga_signals.g0_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_x2_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110011001"
        )
    port map (
            in0 => \N__33127\,
            in1 => \N__33002\,
            in2 => \_gnd_net_\,
            in3 => \N__32934\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_10_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_0_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001000000"
        )
    port map (
            in0 => \N__29954\,
            in1 => \N__33408\,
            in2 => \N__29948\,
            in3 => \N__33611\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_6_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__29945\,
            in1 => \N__29933\,
            in2 => \N__29927\,
            in3 => \N__32891\,
            lcout => \this_vga_signals.g0_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_7_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__29924\,
            in1 => \N__29918\,
            in2 => \N__30149\,
            in3 => \N__29981\,
            lcout => \this_vga_signals.if_N_10_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_7_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101000010"
        )
    port map (
            in0 => \N__31528\,
            in1 => \N__30565\,
            in2 => \N__30487\,
            in3 => \N__31664\,
            lcout => \this_vga_signals.g0_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_o2_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100101011"
        )
    port map (
            in0 => \N__31666\,
            in1 => \N__33877\,
            in2 => \N__31422\,
            in3 => \N__30282\,
            lcout => \this_vga_signals.mult1_un61_sum_c2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010000101011"
        )
    port map (
            in0 => \N__31527\,
            in1 => \N__30564\,
            in2 => \N__30486\,
            in3 => \N__31663\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_N_3L3_1_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100010"
        )
    port map (
            in0 => \N__29900\,
            in1 => \N__31751\,
            in2 => \N__29894\,
            in3 => \N__30182\,
            lcout => \this_vga_signals.g0_41_N_3L3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x0_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101100110011"
        )
    port map (
            in0 => \N__33875\,
            in1 => \N__31526\,
            in2 => \N__33168\,
            in3 => \N__30563\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_c3_x0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_ns_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31037\,
            in2 => \N__30008\,
            in3 => \N__30131\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0,
            ltout => \this_vga_signals_un5_vaddress_if_generate_plus_mult1_un54_sum_c3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_41_N_4L5_1_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001110010"
        )
    port map (
            in0 => \N__33876\,
            in1 => \N__31412\,
            in2 => \N__30005\,
            in3 => \N__31665\,
            lcout => \this_vga_signals.g0_41_N_4L5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \m31_0_x3_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__30281\,
            in1 => \_gnd_net_\,
            in2 => \N__30413\,
            in3 => \_gnd_net_\,
            lcout => \N_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_1_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001111011100"
        )
    port map (
            in0 => \N__30317\,
            in1 => \N__31754\,
            in2 => \N__30635\,
            in3 => \N__30229\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__31409\,
            in1 => \N__31294\,
            in2 => \N__29990\,
            in3 => \N__29987\,
            lcout => \this_vga_signals.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_0_1_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__29975\,
            in1 => \N__30228\,
            in2 => \N__30038\,
            in3 => \N__31753\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_i_o4_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011101000"
        )
    port map (
            in0 => \N__31408\,
            in1 => \N__31293\,
            in2 => \N__29969\,
            in3 => \N__30071\,
            lcout => \this_vga_signals.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_17_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000100000"
        )
    port map (
            in0 => \N__30596\,
            in1 => \N__30399\,
            in2 => \N__31421\,
            in3 => \N__30280\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100001001"
        )
    port map (
            in0 => \N__31145\,
            in1 => \N__33609\,
            in2 => \N__33182\,
            in3 => \N__33411\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_1_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__33931\,
            in1 => \_gnd_net_\,
            in2 => \N__30053\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.g0_0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIE8SF1_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__38267\,
            in1 => \N__34930\,
            in2 => \N__36566\,
            in3 => \N__34993\,
            lcout => \M_last_q_RNIE8SF1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x4_0_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010010110"
        )
    port map (
            in0 => \N__31679\,
            in1 => \N__30509\,
            in2 => \N__30302\,
            in3 => \N__30323\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_5_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_RNIPQ17A7_2_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__31274\,
            in1 => \N__31401\,
            in2 => \N__30050\,
            in3 => \N__30353\,
            lcout => \this_vga_signals.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_6_0_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30026\,
            lcout => \this_vga_signals.g0_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_26_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001101001"
        )
    port map (
            in0 => \N__33415\,
            in1 => \N__34069\,
            in2 => \N__33620\,
            in3 => \N__30602\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_2_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010001000001"
        )
    port map (
            in0 => \N__31130\,
            in1 => \N__33616\,
            in2 => \N__34075\,
            in3 => \N__33414\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2\,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_0_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30020\,
            in3 => \N__33928\,
            lcout => \this_vga_signals.g0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_i_x2_1_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31400\,
            in1 => \N__31273\,
            in2 => \_gnd_net_\,
            in3 => \N__31529\,
            lcout => \this_vga_signals.g0_i_x2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIE5RF1_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36550\,
            in2 => \_gnd_net_\,
            in3 => \N__36104\,
            lcout => \N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_LUT4_0_LC_17_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36933\,
            lcout => \GB_BUFFER_M_this_reset_cond_out_g_0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_3_0_wclke_3_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32209\,
            in1 => \N__32116\,
            in2 => \N__32017\,
            in3 => \N__31911\,
            lcout => \this_spr_ram.mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIO4821_9_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__35267\,
            in1 => \N__33125\,
            in2 => \_gnd_net_\,
            in3 => \N__34649\,
            lcout => \this_vga_signals.m43_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIHT721_6_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__33124\,
            in1 => \N__33926\,
            in2 => \_gnd_net_\,
            in3 => \N__34012\,
            lcout => \this_vga_signals.vaddress_c3_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_5_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110011000110"
        )
    port map (
            in0 => \N__31522\,
            in1 => \N__31678\,
            in2 => \N__30502\,
            in3 => \N__30580\,
            lcout => \this_vga_signals.g0_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIKEN71_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35345\,
            in1 => \N__35253\,
            in2 => \N__34640\,
            in3 => \N__34729\,
            lcout => \this_vga_signals.vaddress_ac0_9_0_a0_1\,
            ltout => \this_vga_signals.vaddress_ac0_9_0_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNI3GK81_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__34831\,
            in1 => \_gnd_net_\,
            in2 => \N__30059\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.CO0_0_i_i\,
            ltout => \this_vga_signals.CO0_0_i_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_a3_0_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001001000"
        )
    port map (
            in0 => \N__32985\,
            in1 => \N__33121\,
            in2 => \N__30056\,
            in3 => \N__32930\,
            lcout => \this_vga_signals.N_7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_RNIL0AS_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__34728\,
            in1 => \N__34622\,
            in2 => \_gnd_net_\,
            in3 => \N__35344\,
            lcout => OPEN,
            ltout => \this_vga_signals.vaddress_c5_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI3GK81_9_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35252\,
            in2 => \N__30161\,
            in3 => \N__34830\,
            lcout => \this_vga_signals.vaddress_9\,
            ltout => \this_vga_signals.vaddress_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_7_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100000100"
        )
    port map (
            in0 => \N__34833\,
            in1 => \N__31064\,
            in2 => \N__30158\,
            in3 => \N__32984\,
            lcout => \this_vga_signals.g1_3_0\,
            ltout => \this_vga_signals.g1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_24_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30155\,
            in3 => \N__33122\,
            lcout => \this_vga_signals.N_7_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_3_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101100000100"
        )
    port map (
            in0 => \N__34832\,
            in1 => \N__31065\,
            in2 => \N__32943\,
            in3 => \N__32986\,
            lcout => \this_vga_signals.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_21_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__31752\,
            in1 => \N__30283\,
            in2 => \_gnd_net_\,
            in3 => \N__31671\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_19_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100000000"
        )
    port map (
            in0 => \N__31407\,
            in1 => \N__30140\,
            in2 => \N__30152\,
            in3 => \N__30167\,
            lcout => \this_vga_signals.mult1_un61_sum_c3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_20_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100110011100"
        )
    port map (
            in0 => \N__31498\,
            in1 => \N__30403\,
            in2 => \N__30498\,
            in3 => \N__30562\,
            lcout => \this_vga_signals.N_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_ns_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33261\,
            in2 => \N__31172\,
            in3 => \N__31178\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_ns\,
            ltout => \this_vga_signals.mult1_un47_sum_axbxc3_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c3_x1_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111010"
        )
    port map (
            in0 => \N__33873\,
            in1 => \N__33079\,
            in2 => \N__30134\,
            in3 => \N__31496\,
            lcout => \this_vga_signals.mult1_un54_sum_c3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_16_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100001001"
        )
    port map (
            in0 => \N__33612\,
            in1 => \N__30689\,
            in2 => \N__33120\,
            in3 => \N__33407\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_c2_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101010111011"
        )
    port map (
            in0 => \N__33874\,
            in1 => \N__31033\,
            in2 => \N__33149\,
            in3 => \N__30560\,
            lcout => \this_vga_signals.mult1_un54_sum_c2_0\,
            ltout => \this_vga_signals.mult1_un54_sum_c2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_40_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__30561\,
            in1 => \_gnd_net_\,
            in2 => \N__30188\,
            in3 => \N__31497\,
            lcout => \this_vga_signals.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_1_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31719\,
            in2 => \_gnd_net_\,
            in3 => \N__31662\,
            lcout => OPEN,
            ltout => \this_vga_signals.g1_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_34_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000100000"
        )
    port map (
            in0 => \N__31411\,
            in1 => \N__30393\,
            in2 => \N__30185\,
            in3 => \N__30276\,
            lcout => \this_vga_signals.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_5_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31718\,
            in2 => \_gnd_net_\,
            in3 => \N__31660\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_38_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000100000"
        )
    port map (
            in0 => \N__31410\,
            in1 => \N__30392\,
            in2 => \N__30176\,
            in3 => \N__30275\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_ns_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31043\,
            in1 => \N__31076\,
            in2 => \_gnd_net_\,
            in3 => \N__30557\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_0_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100010101"
        )
    port map (
            in0 => \N__31720\,
            in1 => \N__30173\,
            in2 => \N__30338\,
            in3 => \N__30227\,
            lcout => \this_vga_signals.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_5_N_2L1_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101111010100"
        )
    port map (
            in0 => \N__31499\,
            in1 => \N__30559\,
            in2 => \N__30503\,
            in3 => \N__31661\,
            lcout => \this_vga_signals.g0_5_5_N_2L1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__33595\,
            in2 => \N__33927\,
            in3 => \N__31793\,
            lcout => this_vga_signals_un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_3_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010001000001"
        )
    port map (
            in0 => \N__31129\,
            in1 => \N__33614\,
            in2 => \N__34076\,
            in3 => \N__33412\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_1_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31736\,
            in2 => \_gnd_net_\,
            in3 => \N__31677\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_28_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001000000"
        )
    port map (
            in0 => \N__30279\,
            in1 => \N__31426\,
            in2 => \N__30326\,
            in3 => \N__30398\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_39_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001000000"
        )
    port map (
            in0 => \N__30397\,
            in1 => \N__31604\,
            in2 => \N__31427\,
            in3 => \N__30278\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_d_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_4_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__31737\,
            in1 => \N__31807\,
            in2 => \N__30311\,
            in3 => \N__30221\,
            lcout => \this_vga_signals.g0_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_5_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30220\,
            in1 => \N__30293\,
            in2 => \N__30412\,
            in3 => \N__30277\,
            lcout => \this_vga_signals.g0_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_0_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101010001"
        )
    port map (
            in0 => \N__31735\,
            in1 => \N__30236\,
            in2 => \N__31808\,
            in3 => \N__30219\,
            lcout => OPEN,
            ltout => \this_vga_signals.g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_4_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110011010"
        )
    port map (
            in0 => \N__30665\,
            in1 => \N__30656\,
            in2 => \N__30650\,
            in3 => \N__31676\,
            lcout => \this_vga_signals.N_5_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_1_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31524\,
            in1 => \N__31289\,
            in2 => \_gnd_net_\,
            in3 => \N__30582\,
            lcout => \this_vga_signals.g0_29_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_22_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010001000001"
        )
    port map (
            in0 => \N__30647\,
            in1 => \N__33615\,
            in2 => \N__34074\,
            in3 => \N__33416\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33930\,
            in2 => \N__30638\,
            in3 => \N__32252\,
            lcout => \this_vga_signals.g3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_33_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30619\,
            lcout => \this_vga_signals.N_7_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_1_2_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__31721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31675\,
            lcout => \this_vga_signals.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_1_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__31525\,
            in1 => \N__30499\,
            in2 => \_gnd_net_\,
            in3 => \N__30583\,
            lcout => \this_vga_signals.g1_0\,
            ltout => \this_vga_signals.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_29_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__30500\,
            in1 => \N__30428\,
            in2 => \N__30422\,
            in3 => \N__30418\,
            lcout => \this_vga_signals.g0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_7_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30347\,
            lcout => \this_reset_cond.M_stage_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_9_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30800\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \M_this_reset_cond_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_reset_cond.M_stage_q_8_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__30799\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30734\,
            lcout => \this_reset_cond.M_stage_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39369\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_2_0_wclke_3_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__32217\,
            in1 => \N__31912\,
            in2 => \N__32031\,
            in3 => \N__32117\,
            lcout => \this_spr_ram.mem_WE_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_4_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39322\,
            ce => \N__34491\,
            sr => \N__34428\
        );

    \this_vga_signals.M_vcounter_q_esr_6_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34539\,
            lcout => \this_vga_signals_M_vcounter_q_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39322\,
            ce => \N__34491\,
            sr => \N__34428\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_5_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31572\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39322\,
            ce => \N__34491\,
            sr => \N__34428\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_7_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110011100"
        )
    port map (
            in0 => \N__34837\,
            in1 => \N__31082\,
            in2 => \N__31070\,
            in3 => \N__32942\,
            lcout => \this_vga_signals.N_12_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIF1T_4_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30683\,
            in3 => \N__30674\,
            lcout => \this_vga_signals.vaddress_c2\,
            ltout => \this_vga_signals.vaddress_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_7_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__34626\,
            in1 => \N__33980\,
            in2 => \N__30668\,
            in3 => \N__34730\,
            lcout => \this_vga_signals.vaddress_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_27_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001000100001"
        )
    port map (
            in0 => \N__33613\,
            in1 => \N__31122\,
            in2 => \N__34017\,
            in3 => \N__33384\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_5_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__31103\,
            in1 => \_gnd_net_\,
            in2 => \N__31097\,
            in3 => \N__33939\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0_6_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__35184\,
            in1 => \N__35313\,
            in2 => \N__32861\,
            in3 => \N__32882\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1_9_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__35312\,
            in1 => \N__32856\,
            in2 => \_gnd_net_\,
            in3 => \N__35183\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNI1TB1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNI65531_0_7_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110110"
        )
    port map (
            in0 => \N__34731\,
            in1 => \N__34627\,
            in2 => \N__34016\,
            in3 => \N__34836\,
            lcout => \this_vga_signals.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x0_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010011011011"
        )
    port map (
            in0 => \N__33479\,
            in1 => \N__33440\,
            in2 => \N__33254\,
            in3 => \N__31781\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g1_5_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010010010"
        )
    port map (
            in0 => \N__32983\,
            in1 => \N__32929\,
            in2 => \N__31069\,
            in3 => \N__34835\,
            lcout => \this_vga_signals.g1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc3_1_x1_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__33478\,
            in1 => \N__33442\,
            in2 => \N__33253\,
            in3 => \N__31782\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc3_1_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001011010"
        )
    port map (
            in0 => \N__31783\,
            in1 => \N__33238\,
            in2 => \N__31598\,
            in3 => \N__33295\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc1_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__33237\,
            in1 => \N__33474\,
            in2 => \_gnd_net_\,
            in3 => \N__33441\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34_6_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31451\,
            in1 => \N__31445\,
            in2 => \_gnd_net_\,
            in3 => \N__34834\,
            lcout => OPEN,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNIQD34Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1_6_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001100110"
        )
    port map (
            in0 => \N__33532\,
            in1 => \N__33473\,
            in2 => \N__31439\,
            in3 => \N__32831\,
            lcout => \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6\,
            ltout => \this_vga_signals.M_vcounter_q_fast_esr_RNIN1DJ1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x0_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101101001"
        )
    port map (
            in0 => \N__31594\,
            in1 => \N__33901\,
            in2 => \N__31436\,
            in3 => \N__33294\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_42_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010110100110"
        )
    port map (
            in0 => \N__31433\,
            in1 => \N__31399\,
            in2 => \N__31295\,
            in3 => \N__31193\,
            lcout => \this_vga_signals.N_5786_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x0_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010110"
        )
    port map (
            in0 => \N__33475\,
            in1 => \N__33358\,
            in2 => \N__33573\,
            in3 => \N__33292\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_x0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un47_sum_axbxc3_x1_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__33356\,
            in2 => \N__33572\,
            in3 => \N__33476\,
            lcout => \this_vga_signals.mult1_un47_sum_axbxc3_x1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIC5EK3_0_7_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110011001"
        )
    port map (
            in0 => \N__31163\,
            in1 => \N__33001\,
            in2 => \_gnd_net_\,
            in3 => \N__32944\,
            lcout => \this_vga_signals.N_12_0\,
            ltout => \this_vga_signals.N_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_ac0_3_c_0_1_0_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000100101"
        )
    port map (
            in0 => \N__33536\,
            in1 => \N__33357\,
            in2 => \N__31133\,
            in3 => \N__33083\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un61_sum_axb1_0_1_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000110001110"
        )
    port map (
            in0 => \N__33477\,
            in1 => \N__33443\,
            in2 => \N__33266\,
            in3 => \N__33359\,
            lcout => \this_vga_signals.mult1_un61_sum_axb1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_5_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31573\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39345\,
            ce => \N__34509\,
            sr => \N__34430\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_x1_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__31593\,
            in1 => \N__31787\,
            in2 => \N__33943\,
            in3 => \N__33296\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc1_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axbxc1_ns_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33265\,
            in1 => \_gnd_net_\,
            in2 => \N__31766\,
            in3 => \N__31763\,
            lcout => \this_vga_signals.mult1_un54_sum_axbxc1_ns\,
            ltout => \this_vga_signals.mult1_un54_sum_axbxc1_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_2_2_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31682\,
            in3 => \N__31667\,
            lcout => \this_vga_signals.g0_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un54_sum_axb1_s_0_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33640\,
            in2 => \_gnd_net_\,
            in3 => \N__33659\,
            lcout => \this_vga_signals.mult1_un54_sum_axb1_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31577\,
            lcout => \this_vga_signals.M_vcounter_q_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39354\,
            ce => \N__34510\,
            sr => \N__34432\
        );

    \this_start_data_delay.M_last_q_RNI1KH61_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__31550\,
            in1 => \N__35539\,
            in2 => \N__33701\,
            in3 => \N__36616\,
            lcout => \this_start_data_delay.N_380\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_d_0_sqmuxa_2_0_a4_0_a2_0_a2_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__34327\,
            in1 => \N__34350\,
            in2 => \N__33776\,
            in3 => \N__34367\,
            lcout => OPEN,
            ltout => \M_this_state_d_0_sqmuxa_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_substate_q_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__34368\,
            in1 => \N__38007\,
            in2 => \N__32300\,
            in3 => \N__35921\,
            lcout => \M_this_substate_qZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39362\,
            ce => 'H',
            sr => \N__36812\
        );

    \this_start_data_delay.M_last_q_RNIO2A13_0_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__36617\,
            in1 => \N__38334\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_233_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIHUID5_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__35909\,
            in1 => \N__37045\,
            in2 => \N__32297\,
            in3 => \N__36935\,
            lcout => \N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_23_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000000110"
        )
    port map (
            in0 => \N__33594\,
            in1 => \N__32264\,
            in2 => \N__33131\,
            in3 => \N__33413\,
            lcout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICPQ11_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36565\,
            in2 => \_gnd_net_\,
            in3 => \N__36134\,
            lcout => \N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_1_3_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35469\,
            lcout => \this_start_data_delay.N_467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_4_0_wclke_3_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__32205\,
            in1 => \N__32103\,
            in2 => \N__32016\,
            in3 => \N__31918\,
            lcout => \this_spr_ram.mem_WE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_spr_ram.mem_mem_5_0_wclke_3_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__32177\,
            in1 => \N__32081\,
            in2 => \N__31996\,
            in3 => \N__31913\,
            lcout => \this_spr_ram.mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIPTJA2_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__37891\,
            in1 => \N__35131\,
            in2 => \N__38737\,
            in3 => \N__38278\,
            lcout => \M_this_spr_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_ppu.oam_cache.read_data_RNI5QFJ1_1_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32735\,
            in1 => \N__32723\,
            in2 => \_gnd_net_\,
            in3 => \N__32693\,
            lcout => \M_this_ppu_spr_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_0_12_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38348\,
            in2 => \_gnd_net_\,
            in3 => \N__35712\,
            lcout => \this_start_data_delay.N_284_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNILPJA2_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__37766\,
            in1 => \N__35130\,
            in2 => \N__38896\,
            in3 => \N__38281\,
            lcout => \M_this_spr_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_6_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001111"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__32879\,
            in2 => \N__32860\,
            in3 => \N__35306\,
            lcout => \this_vga_signals.m47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_6_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34546\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39337\,
            ce => \N__34498\,
            sr => \N__34429\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_9_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34564\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39337\,
            ce => \N__34498\,
            sr => \N__34429\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_7_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34771\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39337\,
            ce => \N__34498\,
            sr => \N__34429\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_8_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34672\,
            lcout => \this_vga_signals.M_vcounter_q_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39337\,
            ce => \N__34498\,
            sr => \N__34429\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_1_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001100"
        )
    port map (
            in0 => \N__32880\,
            in1 => \N__32854\,
            in2 => \N__35189\,
            in3 => \N__35314\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_0_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011111110101"
        )
    port map (
            in0 => \N__35230\,
            in1 => \N__34828\,
            in2 => \N__33272\,
            in3 => \N__35307\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un40_sum_ac0_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011010000"
        )
    port map (
            in0 => \N__34829\,
            in1 => \N__34628\,
            in2 => \N__33269\,
            in3 => \N__35150\,
            lcout => \this_vga_signals.mult1_un40_sum_c3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_30_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000011010"
        )
    port map (
            in0 => \N__33194\,
            in1 => \N__33380\,
            in2 => \N__33582\,
            in3 => \N__33078\,
            lcout => OPEN,
            ltout => \this_vga_signals.mult1_un61_sum_ac0_3_c_0_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIE9FPA_4_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33903\,
            in2 => \N__33212\,
            in3 => \N__33008\,
            lcout => \this_vga_signals.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_35_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33077\,
            lcout => OPEN,
            ltout => \this_vga_signals.N_7_1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_RNIOLNC5_6_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000001001"
        )
    port map (
            in0 => \N__34019\,
            in1 => \N__33546\,
            in2 => \N__33011\,
            in3 => \N__33370\,
            lcout => \this_vga_signals.G_5_i_o2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_32_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000101000"
        )
    port map (
            in0 => \N__33782\,
            in1 => \N__32996\,
            in2 => \N__34784\,
            in3 => \N__32948\,
            lcout => \this_vga_signals.N_19_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIAFQ1_1_6_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001000101"
        )
    port map (
            in0 => \N__32881\,
            in1 => \N__32855\,
            in2 => \N__35315\,
            in3 => \N__35181\,
            lcout => OPEN,
            ltout => \this_vga_signals.m47_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_fast_esr_RNIDJ05_7_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110010001100"
        )
    port map (
            in0 => \N__35182\,
            in1 => \N__32830\,
            in2 => \N__34079\,
            in3 => \N__34827\,
            lcout => \this_vga_signals.SUM_2\,
            ltout => \this_vga_signals.SUM_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_a7_1_3_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000100"
        )
    port map (
            in0 => \N__34018\,
            in1 => \N__33902\,
            in2 => \N__33785\,
            in3 => \N__33545\,
            lcout => \this_vga_signals.g0_0_i_a7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d28_0_a2_0_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33719\,
            in1 => \N__33764\,
            in2 => \N__33746\,
            in3 => \N__35540\,
            lcout => \N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1_6_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__33763\,
            in1 => \N__33742\,
            in2 => \_gnd_net_\,
            in3 => \N__33718\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIHKHB_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33635\,
            in2 => \_gnd_net_\,
            in3 => \N__33657\,
            lcout => \this_vga_signals.vaddress_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_4_rep1_esr_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33689\,
            lcout => \this_vga_signals.M_vcounter_q_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39355\,
            ce => \N__34511\,
            sr => \N__34433\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNIBS0H_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__35342\,
            in1 => \N__33636\,
            in2 => \_gnd_net_\,
            in3 => \N__33656\,
            lcout => \this_vga_signals.vaddress_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_5_rep1_esr_RNI88ES_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010011"
        )
    port map (
            in0 => \N__33658\,
            in1 => \N__34733\,
            in2 => \N__33641\,
            in3 => \N__35343\,
            lcout => \this_vga_signals.vaddress_7\,
            ltout => \this_vga_signals.vaddress_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_m2_0_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011001100000"
        )
    port map (
            in0 => \N__33472\,
            in1 => \N__33439\,
            in2 => \N__33419\,
            in3 => \N__33355\,
            lcout => \this_vga_signals.if_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIK6R81_0_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35607\,
            in1 => \N__38229\,
            in2 => \_gnd_net_\,
            in3 => \N__36562\,
            lcout => \this_start_data_delay.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIGR6G1_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__36563\,
            in1 => \N__36953\,
            in2 => \N__36035\,
            in3 => \N__37997\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_345_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_1_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__35417\,
            in1 => \N__35476\,
            in2 => \N__34100\,
            in3 => \N__35363\,
            lcout => \M_this_state_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIH1242_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__36952\,
            in1 => \N__36564\,
            in2 => \N__35713\,
            in3 => \N__36632\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_12_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__34097\,
            in1 => \N__36166\,
            in2 => \N__34088\,
            in3 => \N__34903\,
            lcout => \M_this_state_qZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39363\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_6_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__34301\,
            in1 => \N__35963\,
            in2 => \N__34379\,
            in3 => \N__36165\,
            lcout => \M_this_state_qZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINO621_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36568\,
            in2 => \_gnd_net_\,
            in3 => \N__36937\,
            lcout => \this_start_data_delay.N_23_1_0\,
            ltout => \this_start_data_delay.N_23_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIMS691_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34085\,
            in3 => \N__36086\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_3_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__34352\,
            in1 => \N__34370\,
            in2 => \N__34082\,
            in3 => \N__35366\,
            lcout => \M_this_state_qZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1_6_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__36938\,
            in1 => \N__34326\,
            in2 => \N__35507\,
            in3 => \N__37979\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_0_i_0_i_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIGTHM1_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__37978\,
            in1 => \N__34299\,
            in2 => \N__34328\,
            in3 => \N__36939\,
            lcout => \this_start_data_delay.N_386\,
            ltout => \this_start_data_delay.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_2_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__34369\,
            in1 => \N__34351\,
            in2 => \N__34331\,
            in3 => \N__34289\,
            lcout => \M_this_state_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39370\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOVDB1_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011000100"
        )
    port map (
            in0 => \N__34325\,
            in1 => \N__34300\,
            in2 => \N__35424\,
            in3 => \N__35459\,
            lcout => \N_465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNILR691_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35961\,
            in2 => \_gnd_net_\,
            in3 => \N__36055\,
            lcout => \this_start_data_delay.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNINRJA2_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__37651\,
            in1 => \N__35135\,
            in2 => \N__37331\,
            in3 => \N__38279\,
            lcout => \M_this_spr_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_0_a2_0_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__35726\,
            in1 => \N__36593\,
            in2 => \N__34916\,
            in3 => \N__35660\,
            lcout => OPEN,
            ltout => \dma_axb0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dma_c4_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__34850\,
            in1 => \N__34940\,
            in2 => \N__34181\,
            in3 => \N__34106\,
            lcout => dma_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_3_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__35611\,
            in1 => \N__38280\,
            in2 => \_gnd_net_\,
            in3 => \N__35144\,
            lcout => dma_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_g0_0_i_o2_0_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__35239\,
            in1 => \N__34716\,
            in2 => \N__34632\,
            in3 => \N__34841\,
            lcout => \this_vga_signals.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_vcounter_q_esr_7_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34775\,
            lcout => \this_vga_signals_M_vcounter_q_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39346\,
            ce => \N__34508\,
            sr => \N__34431\
        );

    \this_vga_signals.M_vcounter_q_esr_8_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34676\,
            lcout => \this_vga_signals_M_vcounter_q_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39346\,
            ce => \N__34508\,
            sr => \N__34431\
        );

    \this_vga_signals.M_vcounter_q_esr_9_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34568\,
            lcout => \this_vga_signals.M_vcounter_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39346\,
            ce => \N__34508\,
            sr => \N__34431\
        );

    \this_vga_signals.M_vcounter_q_6_rep1_esr_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34547\,
            lcout => \this_vga_signals.M_vcounter_q_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39346\,
            ce => \N__34508\,
            sr => \N__34431\
        );

    \M_this_state_q_13_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__35972\,
            in1 => \N__34892\,
            in2 => \N__36992\,
            in3 => \N__35714\,
            lcout => \M_this_state_qZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_11_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__35971\,
            in1 => \N__36421\,
            in2 => \N__36991\,
            in3 => \N__34984\,
            lcout => \M_this_state_qZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39356\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_6__m6_i_a4_0_a2_2_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38285\,
            lcout => OPEN,
            ltout => \N_422_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_6__N_458_i_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__34893\,
            in1 => \N__34985\,
            in2 => \N__34403\,
            in3 => \N__37939\,
            lcout => \N_458_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.un5_vaddress_if_generate_plus_mult1_un40_sum_ac0_3_1_1_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010111"
        )
    port map (
            in0 => \N__35336\,
            in1 => \N__35311\,
            in2 => \N__35251\,
            in3 => \N__35185\,
            lcout => \this_vga_signals.mult1_un40_sum_ac0_3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_i_0_o4_10_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__34974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36130\,
            lcout => \this_start_data_delay.N_242_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_1_3_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35695\,
            in1 => \N__34973\,
            in2 => \N__34894\,
            in3 => \N__36413\,
            lcout => \this_start_data_delay.un20_i_a4_0_a2_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_i_0_a2_2_4_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__35480\,
            in1 => \N__35425\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.N_387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIJNJA2_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__38116\,
            in1 => \N__35120\,
            in2 => \N__37521\,
            in3 => \N__38284\,
            lcout => \M_this_spr_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_0_o2_1_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36414\,
            in2 => \_gnd_net_\,
            in3 => \N__35652\,
            lcout => \this_start_data_delay.N_245_0\,
            ltout => \this_start_data_delay.N_245_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_0_a2_1_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__36161\,
            in1 => \N__34986\,
            in2 => \N__34943\,
            in3 => \N__35983\,
            lcout => un20_i_a4_0_a2_0_a2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_2_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35710\,
            in1 => \N__36097\,
            in2 => \N__34907\,
            in3 => \N__35653\,
            lcout => un20_i_a4_0_a2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNICVMT3_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__35654\,
            in1 => \N__36631\,
            in2 => \N__38141\,
            in3 => \N__36954\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_srsts_i_i_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_7_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__35805\,
            in1 => \N__38228\,
            in2 => \N__35729\,
            in3 => \N__35655\,
            lcout => \M_this_state_qZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_0_a2_2_0_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__38227\,
            in1 => \N__36007\,
            in2 => \_gnd_net_\,
            in3 => \N__36085\,
            lcout => \this_start_data_delay.un20_i_a4_0_a2_0_a2_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_data_count_qlde_i_o4_0_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__35711\,
            in1 => \_gnd_net_\,
            in2 => \N__35669\,
            in3 => \_gnd_net_\,
            lcout => \this_start_data_delay.N_246_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_8_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__35656\,
            in1 => \N__35965\,
            in2 => \N__36984\,
            in3 => \N__35620\,
            lcout => \M_this_state_qZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_vga_signals.M_this_state_d28_0_a2_0_1_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35558\,
            lcout => \this_vga_signals_M_this_state_d28_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_RNIKV6G1_2_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__36936\,
            in1 => \N__36084\,
            in2 => \N__36572\,
            in3 => \N__36054\,
            lcout => \N_1264_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_4_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__38160\,
            in1 => \N__35365\,
            in2 => \N__35503\,
            in3 => \N__35964\,
            lcout => \M_this_state_qZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIOU691_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35962\,
            in2 => \_gnd_net_\,
            in3 => \N__36126\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_337_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_5_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__35460\,
            in1 => \N__35413\,
            in2 => \N__35369\,
            in3 => \N__35364\,
            lcout => \M_this_state_qZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39377\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_ext_address_d_0_sqmuxa_1_0_a4_0_o2_i_o4_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36160\,
            in1 => \N__38159\,
            in2 => \_gnd_net_\,
            in3 => \N__36125\,
            lcout => \this_start_data_delay.N_239_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.un20_i_a4_0_a2_3_0_a4_1_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36083\,
            in2 => \_gnd_net_\,
            in3 => \N__36053\,
            lcout => \this_start_data_delay.N_420_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36020\,
            in2 => \_gnd_net_\,
            in3 => \N__35984\,
            lcout => \N_466\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIVPN44_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__38344\,
            in1 => \N__35904\,
            in2 => \N__37996\,
            in3 => \N__35960\,
            lcout => OPEN,
            ltout => \this_start_data_delay.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_0_LC_21_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__35885\,
            in1 => \N__37983\,
            in2 => \N__35924\,
            in3 => \N__35920\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1_0_0_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__38345\,
            in1 => \N__35905\,
            in2 => \N__37938\,
            in3 => \N__36950\,
            lcout => \this_start_data_delay.M_this_state_q_srsts_0_0_0_a2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_ext_address_q_0_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37090\,
            in1 => \N__35851\,
            in2 => \N__35879\,
            in3 => \N__35878\,
            lcout => \M_this_ext_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_21_24_0_\,
            carryout => \un1_M_this_ext_address_q_cry_0\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_1_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37094\,
            in1 => \N__35827\,
            in2 => \_gnd_net_\,
            in3 => \N__35816\,
            lcout => \M_this_ext_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_0\,
            carryout => \un1_M_this_ext_address_q_cry_1\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_2_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37091\,
            in1 => \N__36382\,
            in2 => \_gnd_net_\,
            in3 => \N__36371\,
            lcout => \M_this_ext_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_1\,
            carryout => \un1_M_this_ext_address_q_cry_2\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_3_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37095\,
            in1 => \N__36355\,
            in2 => \_gnd_net_\,
            in3 => \N__36344\,
            lcout => \M_this_ext_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_2\,
            carryout => \un1_M_this_ext_address_q_cry_3\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_4_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37092\,
            in1 => \N__36328\,
            in2 => \_gnd_net_\,
            in3 => \N__36317\,
            lcout => \M_this_ext_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_3\,
            carryout => \un1_M_this_ext_address_q_cry_4\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_5_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37096\,
            in1 => \N__36301\,
            in2 => \_gnd_net_\,
            in3 => \N__36290\,
            lcout => \M_this_ext_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_4\,
            carryout => \un1_M_this_ext_address_q_cry_5\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_6_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37093\,
            in1 => \N__36271\,
            in2 => \_gnd_net_\,
            in3 => \N__36260\,
            lcout => \M_this_ext_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_5\,
            carryout => \un1_M_this_ext_address_q_cry_6\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_7_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37097\,
            in1 => \N__36241\,
            in2 => \_gnd_net_\,
            in3 => \N__36230\,
            lcout => \M_this_ext_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_6\,
            carryout => \un1_M_this_ext_address_q_cry_7\,
            clk => \N__39397\,
            ce => 'H',
            sr => \N__36815\
        );

    \M_this_ext_address_q_8_LC_21_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__38117\,
            in1 => \N__37082\,
            in2 => \N__36217\,
            in3 => \N__36200\,
            lcout => \M_this_ext_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_21_25_0_\,
            carryout => \un1_M_this_ext_address_q_cry_8\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_9_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37751\,
            in1 => \N__37086\,
            in2 => \N__36190\,
            in3 => \N__36173\,
            lcout => \M_this_ext_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_8\,
            carryout => \un1_M_this_ext_address_q_cry_9\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_10_LC_21_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37632\,
            in1 => \N__37083\,
            in2 => \N__37243\,
            in3 => \N__37226\,
            lcout => \M_this_ext_address_qZ0Z_10\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_9\,
            carryout => \un1_M_this_ext_address_q_cry_10\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_11_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37874\,
            in1 => \N__37087\,
            in2 => \N__37210\,
            in3 => \N__37193\,
            lcout => \M_this_ext_address_qZ0Z_11\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_10\,
            carryout => \un1_M_this_ext_address_q_cry_11\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_12_LC_21_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37499\,
            in1 => \N__37084\,
            in2 => \N__37180\,
            in3 => \N__37163\,
            lcout => \M_this_ext_address_qZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_11\,
            carryout => \un1_M_this_ext_address_q_cry_12\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_13_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__38903\,
            in1 => \N__37088\,
            in2 => \N__37150\,
            in3 => \N__37133\,
            lcout => \M_this_ext_address_qZ0Z_13\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_12\,
            carryout => \un1_M_this_ext_address_q_cry_13\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_14_LC_21_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__37340\,
            in1 => \N__37085\,
            in2 => \N__37117\,
            in3 => \N__37100\,
            lcout => \M_this_ext_address_qZ0Z_14\,
            ltout => OPEN,
            carryin => \un1_M_this_ext_address_q_cry_13\,
            carryout => \un1_M_this_ext_address_q_cry_14\,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \M_this_ext_address_q_15_LC_21_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__37003\,
            in1 => \N__37089\,
            in2 => \N__38773\,
            in3 => \N__37022\,
            lcout => \M_this_ext_address_qZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39403\,
            ce => 'H',
            sr => \N__36818\
        );

    \this_start_data_delay.M_last_q_RNIO2A13_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__36629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38346\,
            lcout => \this_start_data_delay.N_231_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIJ68N1_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__36951\,
            in1 => \N__36591\,
            in2 => \N__36422\,
            in3 => \N__36630\,
            lcout => OPEN,
            ltout => \this_start_data_delay.M_this_state_q_srsts_i_i_0_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_state_q_10_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000000100000"
        )
    port map (
            in0 => \N__36592\,
            in1 => \N__38347\,
            in2 => \N__36575\,
            in3 => \N__36543\,
            lcout => \M_this_state_qZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_this_state_q_srsts_i_i_a2_1_7_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__38343\,
            in1 => \N__38283\,
            in2 => \_gnd_net_\,
            in3 => \N__38164\,
            lcout => \this_start_data_delay.N_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI497F1_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38127\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38620\,
            lcout => \M_this_map_ram_write_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \led_1_7_6__m7_0_a4_0_a2_0_a2_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38008\,
            in2 => \_gnd_net_\,
            in3 => \N__37943\,
            lcout => led_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI7C7F1_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38624\,
            lcout => \M_this_map_ram_write_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI5A7F1_LC_24_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37752\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38626\,
            lcout => \M_this_map_ram_write_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI6B7F1_LC_24_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37611\,
            lcout => \M_this_map_ram_write_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI8D7F1_LC_24_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37475\,
            lcout => \M_this_map_ram_write_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIAF7F1_LC_24_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37312\,
            lcout => \M_this_map_ram_write_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNI9E7F1_LC_24_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38886\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38618\,
            lcout => \M_this_map_ram_write_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \this_start_data_delay.M_last_q_RNIBG7F1_LC_24_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__38619\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38774\,
            lcout => \M_this_map_ram_write_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \M_this_map_address_q_0_LC_26_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39517\,
            in1 => \N__38509\,
            in2 => \N__38602\,
            in3 => \N__38587\,
            lcout => \M_this_map_address_qZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_26_25_0_\,
            carryout => \un1_M_this_map_address_q_cry_0\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_1_LC_26_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39523\,
            in1 => \N__38479\,
            in2 => \_gnd_net_\,
            in3 => \N__38465\,
            lcout => \M_this_map_address_qZ0Z_1\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_0\,
            carryout => \un1_M_this_map_address_q_cry_1\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_2_LC_26_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39518\,
            in1 => \N__38449\,
            in2 => \_gnd_net_\,
            in3 => \N__38435\,
            lcout => \M_this_map_address_qZ0Z_2\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_1\,
            carryout => \un1_M_this_map_address_q_cry_2\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_3_LC_26_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39524\,
            in1 => \N__38422\,
            in2 => \_gnd_net_\,
            in3 => \N__38408\,
            lcout => \M_this_map_address_qZ0Z_3\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_2\,
            carryout => \un1_M_this_map_address_q_cry_3\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_4_LC_26_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39519\,
            in1 => \N__38392\,
            in2 => \_gnd_net_\,
            in3 => \N__38378\,
            lcout => \M_this_map_address_qZ0Z_4\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_3\,
            carryout => \un1_M_this_map_address_q_cry_4\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_5_LC_26_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39521\,
            in1 => \N__38365\,
            in2 => \_gnd_net_\,
            in3 => \N__38351\,
            lcout => \M_this_map_address_qZ0Z_5\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_4\,
            carryout => \un1_M_this_map_address_q_cry_5\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_6_LC_26_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39520\,
            in1 => \N__39607\,
            in2 => \_gnd_net_\,
            in3 => \N__39593\,
            lcout => \M_this_map_address_qZ0Z_6\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_5\,
            carryout => \un1_M_this_map_address_q_cry_6\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_7_LC_26_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39522\,
            in1 => \N__39577\,
            in2 => \_gnd_net_\,
            in3 => \N__39563\,
            lcout => \M_this_map_address_qZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_M_this_map_address_q_cry_6\,
            carryout => \un1_M_this_map_address_q_cry_7\,
            clk => \N__39424\,
            ce => 'H',
            sr => \N__38956\
        );

    \M_this_map_address_q_8_LC_26_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39525\,
            in1 => \N__39547\,
            in2 => \_gnd_net_\,
            in3 => \N__39533\,
            lcout => \M_this_map_address_qZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_26_26_0_\,
            carryout => \un1_M_this_map_address_q_cry_8\,
            clk => \N__39430\,
            ce => 'H',
            sr => \N__38955\
        );

    \M_this_map_address_q_9_LC_26_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__39448\,
            in1 => \N__39526\,
            in2 => \_gnd_net_\,
            in3 => \N__39464\,
            lcout => \M_this_map_address_qZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__39430\,
            ce => 'H',
            sr => \N__38955\
        );
end \INTERFACE\;
